netcdf _pismsheet_elev_mask {
dimensions:
	time = 1 ;
	x = 76 ;
	y = 141 ;
variables:
	byte mask(time, y, x) ;
		mask:units = "" ;
		mask:coordinates = "lat lon" ;
		mask:flag_meanings = "ice_free_bedrock grounded_ice floating_ice ice_free_ocean" ;
		mask:long_name = "ice-type (ice-free/grounded/floating/ocean) integer mask" ;
		mask:pism_intent = "diagnostic" ;
		mask:flag_values = 0b, 2b, 3b, 4b ;
		mask:grid_mapping = "mapping" ;
	double thk(time, y, x) ;
		thk:units = "m" ;
		thk:valid_min = 0. ;
		thk:coordinates = "lat lon" ;
		thk:long_name = "land ice thickness" ;
		thk:pism_intent = "model_state" ;
		thk:standard_name = "land_ice_thickness" ;
		thk:grid_mapping = "mapping" ;
	double topg(time, y, x) ;
		topg:units = "m" ;
		topg:coordinates = "lat lon" ;
		topg:long_name = "bedrock surface elevation" ;
		topg:pism_intent = "model_state" ;
		topg:standard_name = "bedrock_altitude" ;
		topg:grid_mapping = "mapping" ;
data:

 mask =
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    0, 
    0, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    0, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    0, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    4, 
    0, 
    0, 
    2, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4 ;

 thk =
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    740.32940084779, 
    651.020510093267, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    706.494947091031, 
    778.559402428383, 
    814.116264537032, 
    801.739504676735, 
    990.224207126127, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    977.145382090016, 
    1055.87888920149, 
    895.778394914095, 
    1140.61530224505, 
    727.534616843895, 
    894.815975881069, 
    477.908225931155, 
    568.646788565231, 
    1246.3704694047, 
    924.868731510007, 
    897.64054403342, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    672.091508626054, 
    997.400231074673, 
    1179.12325750035, 
    1296.26418132703, 
    1028.87427217045, 
    604.892541099223, 
    547.628244451089, 
    815.395512012361, 
    785.97421832652, 
    843.245765892873, 
    787.870433240054, 
    745.865457878052, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    516.971241833774, 
    574.929079856995, 
    661.865859686301, 
    815.052405224144, 
    1220.91132491635, 
    965.608342599924, 
    1065.86601865631, 
    884.144654690661, 
    790.238667204518, 
    849.080924037526, 
    564.44687902185, 
    860.987512313408, 
    770.912319748348, 
    769.206277976439, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    676.746277663376, 
    0, 
    544.789465732034, 
    593.270967023791, 
    792.097143328298, 
    898.879029394153, 
    798.943417515091, 
    670.556640188295, 
    1039.26411215906, 
    918.271437860337, 
    723.427044317479, 
    1020.1289738042, 
    1190.18883250059, 
    704.435200572545, 
    840.714877339399, 
    813.132993071006, 
    652.903855852459, 
    866.350961608126, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    701.05591586531, 
    998.687688808512, 
    776.063039869157, 
    516.451554265448, 
    691.586127522817, 
    966.107367055305, 
    1088.24996676222, 
    1043.96720471686, 
    1064.78828663186, 
    1035.86383516999, 
    1283.47603795015, 
    1151.76611505423, 
    1211.42764643721, 
    1587.92428547305, 
    837.188850321479, 
    690.631435376084, 
    896.394803753499, 
    0, 
    661.002437245378, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    814.023587723978, 
    0, 
    527.327692878389, 
    818.675539258469, 
    841.166098851563, 
    970.026094744505, 
    1198.23071927574, 
    1385.08450350585, 
    1157.9859018056, 
    1152.60117276924, 
    1198.29587971017, 
    1232.32905043739, 
    942.185195065032, 
    1295.22299683259, 
    1470.4467986256, 
    1069.3735899934, 
    542.438063447978, 
    666.515239176245, 
    734.530148956401, 
    1079.07422588896, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    769.476634072697, 
    723.055122054427, 
    792.82425522377, 
    710.220334993803, 
    859.32560951443, 
    1200.21032967775, 
    1517.36534371014, 
    1486.24373541519, 
    1363.31161530077, 
    1658.02154056692, 
    1583.73686451238, 
    1560.44007351861, 
    1618.57852424578, 
    1702.88754543045, 
    1599.52510625514, 
    1606.88551129654, 
    1152.06977962778, 
    778.249609517056, 
    730.79727164124, 
    793.173407115827, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    766.110591752444, 
    840.328401982617, 
    900.928741604137, 
    897.915144574975, 
    944.631042102025, 
    1087.51784695879, 
    1395.73948420495, 
    1634.6394401179, 
    1490.13498299992, 
    1291.06089057852, 
    1428.54444143404, 
    1482.83576429753, 
    1555.63185493605, 
    1438.9665399385, 
    1424.2970331137, 
    1386.49537896984, 
    1093.63834525407, 
    1001.61348970081, 
    1078.8332355029, 
    1038.36803342134, 
    1119.51333554626, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    801.46660550228, 
    1014.0015554023, 
    873.226839099915, 
    623.173025604958, 
    914.285977704931, 
    1214.04830934269, 
    1625.75095056823, 
    1692.93432219703, 
    1599.79218583988, 
    1545.04758772811, 
    1728.6654906808, 
    1914.48675866717, 
    1744.30360207369, 
    1689.53874564566, 
    1564.49488238467, 
    1396.33977250241, 
    995.284926778381, 
    690.437572367631, 
    882.98992554823, 
    1045.69152920686, 
    967.96745901725, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    689.792946757798, 
    692.068061489256, 
    757.007786436005, 
    927.157205247509, 
    1100.80608518256, 
    1388.00744413965, 
    1571.61815147037, 
    1644.63913223259, 
    1765.78583239371, 
    1982.90058463521, 
    2037.00625445169, 
    1764.02377085613, 
    1823.35867964923, 
    1614.90196305463, 
    1321.46573010913, 
    1277.17400943817, 
    1216.25667466558, 
    1413.12561598047, 
    1221.06808446444, 
    1173.32616196683, 
    892.942427643247, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    739.810129081766, 
    767.869513903105, 
    793.82451562808, 
    860.178403449483, 
    1169.85432287008, 
    1240.76136057239, 
    1294.01663919259, 
    1512.83694493195, 
    1807.64404619996, 
    1833.64663573387, 
    2049.12416050439, 
    2019.33277948899, 
    1619.23257747613, 
    1699.11077887477, 
    1317.05803959341, 
    1119.75850926573, 
    1442.28343572534, 
    793.555154146578, 
    794.070210809389, 
    896.749768185912, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    645.226359555409, 
    772.291562892813, 
    857.792358100949, 
    1005.32349909195, 
    1324.72258456498, 
    1342.46549703858, 
    1357.52826522705, 
    1569.97880679351, 
    1683.05322806056, 
    1806.43393129379, 
    2202.32979072946, 
    1925.43490014295, 
    1710.08041571785, 
    1415.25485401038, 
    939.82121752843, 
    1076.99532114482, 
    845.351381216885, 
    714.235776008206, 
    691.176533651894, 
    1060.34029796081, 
    756.255577166329, 
    960.144760866256, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    665.914482446004, 
    756.966434586848, 
    836.896310671684, 
    1197.72569300907, 
    1519.6352808972, 
    1711.94843105841, 
    1609.39489128448, 
    1479.54785231383, 
    1769.79021787922, 
    1954.89350328933, 
    2153.32470609964, 
    1703.28145683202, 
    1871.13099869672, 
    1357.50353975343, 
    1182.09637129258, 
    1256.25794156673, 
    1075.71539036336, 
    577.183811545576, 
    1040.03791360855, 
    1076.33865524743, 
    738.582748211793, 
    763.128367216782, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    963.746099283357, 
    583.291536687557, 
    738.149429958358, 
    1085.88300043751, 
    1335.64605432399, 
    1563.12529907415, 
    1657.83091653071, 
    1709.89795912765, 
    1392.16446638156, 
    1767.44391619394, 
    1738.09262725992, 
    2110.39330692384, 
    2052.4199581608, 
    2088.49804489535, 
    1894.88598428794, 
    1821.82666270849, 
    1351.85809874788, 
    1162.85986984937, 
    757.033810822012, 
    880.253679501072, 
    752.55827159958, 
    748.490517245414, 
    953.415184575397, 
    938.069313137424, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    664.185117051632, 
    786.483335606195, 
    699.601241343417, 
    988.766450425168, 
    1380.74819993755, 
    1570.60420451238, 
    1666.00914302491, 
    1663.14675439765, 
    1660.07273358732, 
    1941.8904024516, 
    2056.40733551862, 
    2219.11285481941, 
    2290.40922394733, 
    2276.47427036794, 
    2062.94666574065, 
    1727.4667681731, 
    1538.69776388079, 
    1379.23696962139, 
    1180.12009255133, 
    616.706332048481, 
    826.528041208102, 
    1076.16371712871, 
    595.756512698189, 
    601.476211579043, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    947.30134616487, 
    927.576564953108, 
    777.53467095509, 
    1159.97352553386, 
    1443.95522708837, 
    1540.57488574272, 
    1653.4940934444, 
    1761.98894598281, 
    1903.86557960431, 
    2181.4933209107, 
    2320.32531529931, 
    2348.42806524165, 
    2377.47502821547, 
    2233.76458961367, 
    1993.908155169, 
    1928.32195498921, 
    1795.94955924286, 
    1396.49176302575, 
    1035.38696282088, 
    830.576236196791, 
    608.176944205519, 
    1038.96146319234, 
    1267.50823988534, 
    0, 
    961.431172391549, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    773.504511699971, 
    931.240561392977, 
    914.124033063805, 
    1228.67622453735, 
    1225.0794727404, 
    1485.93671275897, 
    1705.74414637671, 
    1854.71016357165, 
    2003.38057098635, 
    2191.57960726528, 
    2300.62882456309, 
    2295.39178402919, 
    2245.44473394981, 
    2116.11938024876, 
    1940.27703620443, 
    1849.40138598073, 
    2043.61782139474, 
    1534.72219363503, 
    1309.14382385765, 
    1117.80318321462, 
    986.434315444957, 
    961.481921420512, 
    771.089055914368, 
    612.04387195732, 
    1153.77651461266, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    829.342024079655, 
    1036.48922237269, 
    1504.76367376735, 
    1445.60847184085, 
    1593.87039547385, 
    1786.94896627566, 
    1911.41596265927, 
    2016.67181751697, 
    2115.29130667093, 
    2215.32813483864, 
    2247.56720715793, 
    2252.79916598868, 
    2268.62142182312, 
    2135.25124371344, 
    2248.98659010329, 
    2118.94935290094, 
    1656.46370148007, 
    1430.20066345016, 
    1333.86810981001, 
    1330.82149170084, 
    1089.86019624601, 
    1255.78191627885, 
    1339.18545095702, 
    1147.98896915664, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    779.822587598119, 
    910.759907664515, 
    1174.51060254855, 
    1553.48615864834, 
    1507.96957791324, 
    1808.54228001119, 
    1989.53556471927, 
    2074.36826272518, 
    2027.28035490647, 
    2030.8517024486, 
    2120.30102019864, 
    2181.63938364144, 
    2252.10773898076, 
    2391.94951296732, 
    2194.71572818285, 
    1969.53829708238, 
    1847.81885329569, 
    1606.66969939561, 
    1100.53724494336, 
    971.028431787548, 
    1263.49022860995, 
    1343.35818856489, 
    1670.55213076881, 
    1164.49312216302, 
    1166.79620371329, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    853.591929543137, 
    1143.46669943813, 
    1261.69555228853, 
    1240.09521830023, 
    1608.02480215719, 
    1501.41693992614, 
    1865.98753803961, 
    1884.66521796675, 
    1977.6037943205, 
    2080.65974768032, 
    2058.37053544212, 
    2025.46604107451, 
    2047.69297148758, 
    2079.81908395376, 
    2036.54992678912, 
    2039.57065295687, 
    2038.15755624857, 
    1975.99569243522, 
    1677.26336133447, 
    1414.98983182991, 
    1356.86403752403, 
    1401.83660869913, 
    1125.96358816361, 
    690.918333133029, 
    641.063449571816, 
    898.292657705763, 
    696.720792035126, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    789.487757488336, 
    922.188550001941, 
    1204.94896392275, 
    1127.11726894856, 
    1312.98764219661, 
    1160.80110766634, 
    1308.54644227672, 
    1630.68288058746, 
    1669.93248850183, 
    1791.79317770452, 
    2025.00552973435, 
    2013.02598417295, 
    1937.20951132062, 
    1909.93429201636, 
    2038.18176481873, 
    2003.36602516807, 
    2030.17684897352, 
    2025.6624738522, 
    1687.33692517661, 
    1613.46153791905, 
    1524.12406541689, 
    1418.88456537328, 
    1308.03224849181, 
    1235.68198079328, 
    829.832733470305, 
    628.060121278545, 
    885.254330766589, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    731.010447126817, 
    948.705561627144, 
    561.400232190044, 
    1190.47311990612, 
    1367.03271609588, 
    1196.13054886861, 
    923.086896496086, 
    1123.67945236452, 
    1444.67855436406, 
    1542.31766843971, 
    1729.82881988932, 
    1864.82568568936, 
    1994.8430386949, 
    1990.61963046121, 
    1937.54852759429, 
    1949.56728114413, 
    1827.86143362583, 
    1781.63115262315, 
    1913.9205293357, 
    1818.50778485254, 
    1749.21787697488, 
    1459.29938792491, 
    1485.47420887737, 
    1542.9915393325, 
    1099.98755694116, 
    1025.52945517652, 
    1259.42991052772, 
    1141.22552027025, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    762.727179696108, 
    847.066189173929, 
    1186.74576816494, 
    843.146269390191, 
    921.486001572678, 
    1051.11980087088, 
    936.553940297711, 
    1228.84371122646, 
    1496.9993704613, 
    1488.92449965109, 
    1672.76502954809, 
    1904.66435912261, 
    2070.41445195264, 
    2106.5079462957, 
    2070.46732878762, 
    2025.61914538489, 
    1891.66325936628, 
    2008.91050156342, 
    1956.46251039512, 
    1794.39016545806, 
    1977.94367291777, 
    1690.9414722572, 
    1474.1678882353, 
    1352.03691834954, 
    1072.47836991547, 
    1375.8809818216, 
    1403.25708244099, 
    1409.00424525909, 
    1053.35451326569, 
    1155.35217812205, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    529.96246003292, 
    554.482486025395, 
    914.664713980035, 
    987.876730318165, 
    1224.32066100405, 
    1096.4686834232, 
    815.60146887573, 
    1012.09101534968, 
    1329.15008633812, 
    1541.0860901019, 
    1369.68762474992, 
    1538.66106072887, 
    1879.09305919533, 
    2042.3671161265, 
    2119.68813253871, 
    2031.83809140698, 
    1956.79339223939, 
    2008.87881058578, 
    2107.57098294641, 
    1784.05078210003, 
    1960.56899684488, 
    2091.9712027155, 
    1680.49319405285, 
    1522.09586260789, 
    1452.03088359471, 
    1564.56439833697, 
    1406.02824603074, 
    1375.51115138219, 
    1214.44508226583, 
    791.996359112675, 
    994.933776309997, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    723.732454184361, 
    719.365246802671, 
    850.438795207267, 
    576.284144075689, 
    661.273037578639, 
    865.124178217155, 
    1289.37510700975, 
    1564.61615686314, 
    1551.33743839634, 
    1493.76158577699, 
    1744.31873774922, 
    1891.73085874245, 
    2043.66023712329, 
    2102.5111638907, 
    2141.81472335044, 
    2113.44793849684, 
    2053.9761864151, 
    2062.30539260346, 
    2189.09091465333, 
    1891.42424116739, 
    1718.83736939967, 
    1929.16125667894, 
    1884.30170033278, 
    1648.43685700749, 
    1494.21099718014, 
    1391.77221660577, 
    1116.40244659405, 
    734.988611505717, 
    967.357554804067, 
    1107.61101378933, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    699.872051138355, 
    901.336325510045, 
    1282.89279302273, 
    1511.41228842094, 
    1625.35619134769, 
    1652.71168591744, 
    1633.96403131304, 
    1753.4453235198, 
    1769.58479950966, 
    2002.66680139241, 
    2129.77743419275, 
    2138.37366436821, 
    2265.02919862553, 
    2287.5959654266, 
    2274.37918080968, 
    2192.69122045471, 
    2030.57357157477, 
    1841.70132693002, 
    1831.12944161265, 
    1784.80724471083, 
    1756.51440124954, 
    1671.80242899127, 
    1344.30849810349, 
    1144.80842755095, 
    1441.85942286278, 
    1295.25923656503, 
    1156.19279506968, 
    1088.30052926708, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    702.542626939797, 
    736.662387657622, 
    1002.34951779454, 
    1280.40810555484, 
    1479.91197126757, 
    1499.40280033348, 
    1556.39817046852, 
    1559.00980994638, 
    1621.10102219384, 
    1727.46760923562, 
    1990.71991469875, 
    2183.21473240341, 
    2156.576900248, 
    2240.0593533623, 
    2183.69805684058, 
    2229.21717094323, 
    2244.74074155447, 
    2107.28318646292, 
    1896.86172808734, 
    1890.71416148878, 
    1854.15317014889, 
    1829.75516284227, 
    1738.58115766029, 
    1553.56945936068, 
    1457.32232058723, 
    1393.72267516412, 
    968.40560888724, 
    896.740791552496, 
    750.840256998453, 
    842.892305032236, 
    698.646005935741, 
    915.119759085519, 
    852.402875598839, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    674.834103125832, 
    706.674720681005, 
    1021.56813748595, 
    1228.89880005541, 
    1379.71203521524, 
    1491.50120484277, 
    1598.95882063978, 
    1576.75664083018, 
    1584.49399516688, 
    1750.08463307246, 
    1957.73288062655, 
    2107.28548089004, 
    2140.39547092027, 
    2098.49220874292, 
    2025.81102074289, 
    2052.91663444519, 
    2060.33681362602, 
    1939.52204962713, 
    1879.83533944408, 
    1952.20523335271, 
    1943.75012039598, 
    1916.01425582475, 
    1867.03214955368, 
    1712.6824105303, 
    1483.96277881548, 
    1394.45365549702, 
    1073.5755345058, 
    766.94644590151, 
    633.925049988673, 
    1366.84453434019, 
    1211.36021230239, 
    755.568036944489, 
    716.40880969223, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    708.839433120053, 
    788.809076869518, 
    1008.36151513259, 
    1209.04616565599, 
    1376.51721203688, 
    1517.803092067, 
    1683.9633018418, 
    1645.89289242984, 
    1729.82123086183, 
    1767.00595471022, 
    1916.56378490924, 
    2056.69881193472, 
    2125.06059307409, 
    2046.18304451163, 
    2032.132656711, 
    2102.17771564979, 
    2033.80600475594, 
    1926.36196325225, 
    1975.15567838446, 
    2123.17716063684, 
    2009.01435014982, 
    1990.26687270359, 
    2012.58547095171, 
    1921.94757313665, 
    1618.34419067383, 
    1590.94480247395, 
    1396.81478546368, 
    1131.92921598134, 
    910.274830175971, 
    1135.12590692375, 
    1572.95864046019, 
    609.965247037868, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    802.616007798045, 
    769.065155855942, 
    976.72934343125, 
    1244.12159023943, 
    1249.47232541415, 
    1471.2941188809, 
    1602.83468584782, 
    1689.11687742713, 
    1711.03631592933, 
    1843.21354430366, 
    1930.24987996978, 
    2023.08653291242, 
    2213.01049123327, 
    2145.83305283642, 
    2209.83351706356, 
    2185.30573640421, 
    2126.47388977219, 
    2219.8600403561, 
    2105.59991892024, 
    2182.84075786229, 
    2029.55033948969, 
    2200.73275124099, 
    2110.96284296138, 
    1976.95389935017, 
    1848.41107854575, 
    1738.49679040766, 
    1686.26826083464, 
    1478.41443215355, 
    1171.0517444936, 
    1197.48830028105, 
    1771.14543649492, 
    1050.52033079702, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    813.18723375188, 
    1123.02150425706, 
    1167.11280522478, 
    1375.25249195704, 
    1464.83135685302, 
    1589.7547179851, 
    1736.44297165034, 
    1867.49751383098, 
    1950.43374435526, 
    2085.50702900513, 
    2175.30841125978, 
    2245.36966687198, 
    2266.00909809946, 
    2285.79639553963, 
    2304.18788348649, 
    2371.91393297103, 
    2254.87520981262, 
    2267.34879433373, 
    2163.51016281284, 
    2239.84863941808, 
    2134.05844995919, 
    2004.73729130439, 
    2150.65127308277, 
    1824.88610398487, 
    1893.84459472185, 
    1897.36881971494, 
    2055.19058350259, 
    1591.91199171789, 
    994.086367954969, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    703.14005414469, 
    878.273218035964, 
    938.660279717851, 
    1195.99492903569, 
    1306.41983844424, 
    1536.44546354636, 
    1726.62472111012, 
    1845.62091186536, 
    1892.30099101015, 
    2102.51986720419, 
    2192.61901571496, 
    2292.76988115777, 
    2304.59251532883, 
    2283.07666112183, 
    2389.72820134452, 
    2426.16888519213, 
    2420.79598257652, 
    2311.94983508988, 
    2347.59990555756, 
    2245.44739129739, 
    2078.12561302291, 
    2187.8753504493, 
    2239.05431866223, 
    2045.71614583319, 
    2048.33663773911, 
    2037.29271034482, 
    1846.21159760674, 
    1159.05270001727, 
    772.157421911658, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    862.485062942575, 
    997.665754500776, 
    1226.54576074683, 
    1431.89983125685, 
    1689.1704821541, 
    1833.14492496653, 
    1882.0418705423, 
    1916.6138859483, 
    2140.58528609374, 
    2263.0668923903, 
    2317.42431155897, 
    2372.73746651287, 
    2374.9326061699, 
    2473.58912071058, 
    2436.76236018258, 
    2339.65422998288, 
    2432.0347359719, 
    2267.37944061721, 
    2222.78876673016, 
    2292.08659578289, 
    2347.73719511877, 
    2268.02125437662, 
    2151.25679826436, 
    2046.75970623187, 
    1803.25228235223, 
    1303.85723726688, 
    780.447709758619, 
    667.978364342743, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    894.391260020576, 
    1031.35200975023, 
    1300.29075683567, 
    1543.64665435372, 
    1732.51368627545, 
    1829.18773679154, 
    1944.85710703408, 
    2015.74806069272, 
    2083.26345136153, 
    2220.5545933934, 
    2282.83990686878, 
    2336.91294687421, 
    2381.47579702268, 
    2417.44139109817, 
    2269.49261942524, 
    2234.78219457019, 
    2408.23313245633, 
    2364.70431745912, 
    2365.43951053137, 
    2363.05051462206, 
    2454.59700530659, 
    2345.35700600807, 
    2211.48603721666, 
    2052.55593157314, 
    1781.76287461222, 
    1535.35099240584, 
    1278.97427898358, 
    1503.85111958016, 
    461.948379911192, 
    469.799095438841, 
    802.935172419216, 
    973.509729361934, 
    840.36261108746, 
    915.731553087865, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    767.340846726978, 
    947.292256015114, 
    1268.77686051255, 
    1413.68988906867, 
    1575.68360340934, 
    1680.95130886748, 
    1843.13010311743, 
    1919.42996815575, 
    1997.213118908, 
    2122.04458252532, 
    2220.34269357903, 
    2280.10182403339, 
    2287.00714640397, 
    2387.74603550926, 
    2371.8969175851, 
    2426.65253452222, 
    2369.62455640898, 
    2465.46397658031, 
    2466.17132641511, 
    2440.70998526032, 
    2540.08331368613, 
    2508.71970205923, 
    2279.60679754789, 
    2312.19745732958, 
    2069.36310456921, 
    1833.48381828518, 
    1491.60718179202, 
    1133.3468308287, 
    1330.55314363503, 
    1173.553910122, 
    898.016213521143, 
    998.707959630984, 
    534.841689070563, 
    626.671407322524, 
    0, 
    0, 
    1155.82381664277, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    855.262751003474, 
    868.360138742206, 
    1126.64401810743, 
    1308.13739000429, 
    1420.22220566039, 
    1605.42984399971, 
    1678.76188769133, 
    1756.16049658896, 
    1910.85351087235, 
    2009.87172356028, 
    2133.78297678654, 
    2220.29924499212, 
    2261.86555707907, 
    2286.01635839023, 
    2382.8410830684, 
    2368.77324052828, 
    2479.99091909767, 
    2380.05359468491, 
    2484.98646858803, 
    2568.7591752612, 
    2584.34404330385, 
    2595.89607923082, 
    2543.49310279813, 
    2441.09075724097, 
    2300.52708767197, 
    2394.70015788147, 
    2122.88724922013, 
    1673.25048550376, 
    1156.27860566596, 
    1110.08615909237, 
    1141.8227280053, 
    1055.68498403777, 
    1285.58977415245, 
    940.099173954028, 
    636.484203052811, 
    0, 
    0, 
    1074.96585998866, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    837.820448500966, 
    1031.2501599338, 
    1251.45726619613, 
    1351.90309959601, 
    1395.15426577117, 
    1565.93533501521, 
    1637.41377740557, 
    1711.3943410599, 
    1847.06319911482, 
    1993.36534413914, 
    2113.73047293227, 
    2199.33015618605, 
    2221.50435241152, 
    2275.67309826753, 
    2321.80267326564, 
    2366.97857016471, 
    2453.68818649131, 
    2490.76587581206, 
    2560.98577960489, 
    2659.98478797066, 
    2556.11309841336, 
    2527.07445190895, 
    2469.67061951236, 
    2535.93452104413, 
    2610.64107871989, 
    2586.22602578311, 
    2608.16764944869, 
    2153.03567564869, 
    1668.26276536977, 
    1412.24912879483, 
    1386.91856377949, 
    1409.76150934561, 
    1329.66195427639, 
    1000.19965517026, 
    695.535074309979, 
    719.451473177927, 
    837.845111749989, 
    1220.67567062346, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    770.704169178868, 
    818.973009804869, 
    979.619548196021, 
    1253.26018875578, 
    1382.69467452587, 
    1485.88495227564, 
    1598.66007909772, 
    1701.03882664028, 
    1847.02484248881, 
    1982.89893316706, 
    2132.69173297659, 
    2226.37816310341, 
    2209.18973156241, 
    2263.70205590155, 
    2306.91377983127, 
    2361.85487792604, 
    2460.54953061579, 
    2528.05513578309, 
    2491.85272273835, 
    2654.79729874999, 
    2576.06246918841, 
    2511.60358236959, 
    2395.89651734086, 
    2664.72407455952, 
    2785.95418919392, 
    2752.45430845265, 
    2825.78036477596, 
    2405.35168907198, 
    2073.24382504628, 
    1736.88884328618, 
    1682.36159248719, 
    1619.90784712835, 
    1478.50157012658, 
    1603.51400678383, 
    1173.22454940275, 
    851.195227668593, 
    901.213880785241, 
    1127.13018917539, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    674.478564875594, 
    775.651131703533, 
    1080.55905782371, 
    1316.77527951148, 
    1469.66067142899, 
    1570.81873303043, 
    1716.74914363072, 
    1886.31829263459, 
    2100.1131872441, 
    2122.51905011679, 
    2322.99238037393, 
    2196.96254410749, 
    2310.52404015802, 
    2411.18110117478, 
    2441.88858465043, 
    2445.09973336687, 
    2465.79057154706, 
    2635.90441533745, 
    2761.72719725972, 
    2685.08793905466, 
    2630.46240688579, 
    2613.81902244813, 
    2712.62677744483, 
    2768.54274261112, 
    2778.67293265512, 
    2695.82086351822, 
    2486.31072772759, 
    2611.9076826777, 
    2059.6094177189, 
    1744.37838400983, 
    1202.99669349652, 
    1201.00954133498, 
    1490.58202441173, 
    1376.68008121256, 
    855.765807131495, 
    887.635935417921, 
    853.8859841915, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    633.964142849262, 
    787.334513719479, 
    1036.03664402726, 
    1383.44598478046, 
    1603.60752053861, 
    1669.42116150928, 
    1777.42068241016, 
    1877.45842540888, 
    1958.22961796265, 
    2100.70723839082, 
    2241.35961766034, 
    2279.14573599883, 
    2349.71024325289, 
    2497.71777251968, 
    2468.61871207004, 
    2429.70071998259, 
    2519.38492833823, 
    2555.30090327521, 
    2752.37870435488, 
    2744.89392811262, 
    2803.75599846728, 
    2822.08942361554, 
    2855.73639230428, 
    2706.95710103649, 
    2765.60069250747, 
    2532.1002853416, 
    2631.79555729746, 
    2537.59582869376, 
    2224.39903979893, 
    1856.48682361877, 
    1489.16647012251, 
    1264.06440848766, 
    1106.92010219374, 
    882.935328991917, 
    915.854600818732, 
    694.162144670149, 
    0, 
    0, 
    1190.55511290971, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    844.006622235478, 
    875.729384716392, 
    1035.48151513968, 
    1378.00921009952, 
    1612.28235078228, 
    1689.17257871409, 
    1861.20563075652, 
    1867.38865755742, 
    2017.22377869732, 
    2101.41986546489, 
    2206.58396138603, 
    2289.44196832807, 
    2355.38373921478, 
    2457.90575874382, 
    2506.25284428755, 
    2537.28553679981, 
    2607.43716106607, 
    2590.24513735272, 
    2754.04005462542, 
    2729.37135351245, 
    2781.40400962656, 
    2852.00393722846, 
    2997.93926482276, 
    2768.56308336344, 
    2664.92098573923, 
    2619.17918047549, 
    2651.39938336292, 
    2536.72664281452, 
    2353.95997429678, 
    2161.70692508425, 
    2030.93575235362, 
    1681.04618662119, 
    1446.92091929916, 
    1031.87962518696, 
    904.697714993051, 
    821.881571844371, 
    0, 
    0, 
    791.575107716473, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    754.290809794592, 
    935.907589844913, 
    862.000674296646, 
    1119.88537396759, 
    1339.05186582555, 
    1679.89825639866, 
    1856.11788984857, 
    1832.2912797515, 
    1955.46844315604, 
    2109.60657008995, 
    2144.37376572645, 
    2186.28189443705, 
    2275.1390327991, 
    2356.8124656728, 
    2432.73928551176, 
    2569.88090800871, 
    2633.10677125494, 
    2647.94106231832, 
    2618.76895433321, 
    2694.97740508873, 
    2786.45389450115, 
    2876.09713652492, 
    2910.58499043343, 
    2990.23501487103, 
    2825.39707439031, 
    2658.96908202278, 
    2660.76825882433, 
    2800.67103991078, 
    2619.29457133929, 
    2503.95163510348, 
    2220.04509071596, 
    1943.67851721248, 
    1876.53855198578, 
    1488.65453702465, 
    1108.1110165706, 
    900.708422989081, 
    1277.4200799315, 
    585.270334821795, 
    972.409084196659, 
    1389.70368415416, 
    1192.4678680528, 
    971.607389906487, 
    713.48557754912, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    748.103126655991, 
    824.216223822836, 
    901.642410368816, 
    1084.1027943114, 
    1509.477334379, 
    1695.90088537329, 
    1736.18442924934, 
    1872.45564513792, 
    1959.48150070642, 
    2097.21884392533, 
    2129.15079532576, 
    2172.17493774861, 
    2299.16985707071, 
    2393.92073452509, 
    2400.45223500848, 
    2673.63323542618, 
    2719.01259540956, 
    2736.78352802185, 
    2650.16802647748, 
    2552.98777109426, 
    2847.69145621024, 
    2929.04959276222, 
    2949.35297248279, 
    2968.01253873684, 
    2883.32068971197, 
    2855.70286546705, 
    2859.95737100007, 
    2851.88593958971, 
    2733.70899509987, 
    2718.20874573695, 
    2579.41277355035, 
    2693.98869732549, 
    2062.01383972018, 
    1931.86816128941, 
    1539.93069467848, 
    1099.23540806347, 
    1129.2998318215, 
    967.575997186485, 
    1040.33171463585, 
    1748.62328927311, 
    0, 
    0, 
    0, 
    669.187818015947, 
    939.517978408567, 
    743.05989951446, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    626.529976335645, 
    864.623844880338, 
    1012.28753319348, 
    1249.8665286206, 
    1485.81716205772, 
    1579.33094140789, 
    1614.76746726208, 
    1747.88916051814, 
    2010.54477424516, 
    2149.84184340066, 
    2518.56660557035, 
    2278.95991902664, 
    2413.89084541526, 
    2447.08676905922, 
    2504.34567580718, 
    2565.76073169744, 
    2719.16924857105, 
    2803.79147209056, 
    2826.01121788661, 
    2817.19472854943, 
    2848.38187695159, 
    2826.97219691494, 
    2873.16068730802, 
    2897.71223774223, 
    2896.72626767321, 
    2880.56957112712, 
    2873.54276426362, 
    2769.64365867953, 
    2722.51501232624, 
    2780.18955726892, 
    2940.47287145821, 
    2944.00029116348, 
    2290.33365007268, 
    2164.21907661969, 
    1533.50073146507, 
    1197.6920555792, 
    1484.91486720444, 
    1510.50866316341, 
    2003.44252078508, 
    740.303324312754, 
    0, 
    0, 
    641.198580407884, 
    1541.45058157435, 
    1000.78834257153, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    740.931832610591, 
    772.036260075904, 
    993.486596141686, 
    1471.0868521788, 
    1654.46246586912, 
    1592.0075862314, 
    1666.42477918571, 
    1794.55980693706, 
    1932.92849204053, 
    2062.34750242005, 
    2289.21524739603, 
    2409.82839708002, 
    2313.96563175137, 
    2388.43913640482, 
    2503.89957958899, 
    2663.50233304555, 
    2624.56652099189, 
    2694.02801964242, 
    2777.65935167519, 
    2707.93947583723, 
    2669.04422173539, 
    2717.43381712668, 
    2847.14601729271, 
    2813.34018580099, 
    2931.65591077581, 
    2913.3245074284, 
    2822.44151910975, 
    2773.17373985692, 
    2759.5908030825, 
    2814.70840745803, 
    2983.96489508565, 
    2738.67660205286, 
    2101.46120984171, 
    1713.33176683629, 
    1647.19867324929, 
    1915.24185217349, 
    2115.06076781106, 
    2284.43053941499, 
    1377.80868990555, 
    0, 
    0, 
    0, 
    1500.9809036425, 
    1163.73900066436, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    854.606257321113, 
    778.169097675974, 
    988.330277174255, 
    1306.14947532562, 
    1358.67538042818, 
    1703.8826865645, 
    1668.42136224772, 
    2030.39712143721, 
    1884.20951292572, 
    1961.83155351164, 
    2039.60406206901, 
    2202.95702292345, 
    2119.78099861613, 
    2383.48257650118, 
    2521.6115144392, 
    2611.60739039051, 
    2596.83611932913, 
    2736.18176050173, 
    2863.61884559128, 
    2770.18042325942, 
    2825.87406476012, 
    2840.96712110713, 
    2819.48865630996, 
    2837.38028963445, 
    3000.61815115059, 
    2895.83473526022, 
    2831.01367525575, 
    2816.5003216635, 
    2755.4306600559, 
    2744.38654626748, 
    2658.86812079064, 
    2363.25383055864, 
    2027.50714119935, 
    1666.35640818763, 
    1765.90967465499, 
    1945.40014335922, 
    1940.61072125267, 
    2085.72686397927, 
    795.05324292446, 
    0, 
    763.524894275172, 
    625.154787240807, 
    1718.56410727688, 
    751.587821805509, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    829.894308563036, 
    1061.27908969274, 
    1047.26646146725, 
    1282.26164996446, 
    1606.93818046502, 
    1704.09573290597, 
    1773.41270727079, 
    1973.820255025, 
    1979.06089775292, 
    2159.09827042297, 
    2275.66245747398, 
    2345.19970840824, 
    2367.15616963479, 
    2476.35234235321, 
    2601.41362183514, 
    2625.17136459743, 
    2726.43042992347, 
    2842.85900698743, 
    2862.52312943665, 
    2983.84442663978, 
    2952.96096551312, 
    2784.966656576, 
    2944.8283182798, 
    2959.49021791692, 
    2989.85993318238, 
    2939.1920283812, 
    2860.65355291086, 
    2706.28410545386, 
    2656.22758626085, 
    2488.97268063739, 
    2194.00212697417, 
    2305.02914120421, 
    2376.0213407451, 
    2421.11664951336, 
    1909.21690062647, 
    2069.9487004566, 
    1576.71142424545, 
    856.437889381818, 
    705.408895451174, 
    841.044216930187, 
    724.501044408823, 
    1110.35836361617, 
    985.823752387318, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    833.923149261272, 
    1015.25375776309, 
    1013.12507205745, 
    1677.1980587517, 
    1772.15317444728, 
    1736.2972914035, 
    2065.61557237704, 
    1968.1484207722, 
    1967.21698236757, 
    2274.94265119461, 
    2336.12790314334, 
    2433.22438304977, 
    2429.52182776047, 
    2540.72251480537, 
    2705.95697658154, 
    2722.87196281905, 
    2689.38392959796, 
    2765.64593753022, 
    2822.93126506678, 
    2857.28478935912, 
    2898.08217635481, 
    2849.92634346108, 
    2898.26187165082, 
    2964.17391577869, 
    2983.12080049023, 
    2871.0425337345, 
    2854.83576156696, 
    2764.77250963765, 
    2722.74451999628, 
    2549.56934318349, 
    2310.35138076776, 
    2452.92989413179, 
    2308.13777325443, 
    1941.11656818417, 
    1749.51904410475, 
    2017.742643302, 
    1719.65613415446, 
    1403.17931894419, 
    1001.08279199324, 
    790.91675248479, 
    830.615820409138, 
    1006.25251136568, 
    1055.60421079643, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1264.76131382809, 
    1516.65785130975, 
    1635.39206887495, 
    1661.86490953331, 
    1955.67307219291, 
    1972.01055489192, 
    2117.45542454274, 
    2124.56046973083, 
    2261.29551201502, 
    2565.17275380394, 
    2606.01860054326, 
    2605.04961854312, 
    2661.36691084079, 
    2675.6980801795, 
    2663.6368291756, 
    2716.2504067043, 
    2788.07834178724, 
    2788.61023868536, 
    2822.3797280258, 
    2950.78407748392, 
    2936.77913938965, 
    3018.13989669931, 
    2931.87685210448, 
    2915.97240130944, 
    2927.64114994553, 
    2884.53924843412, 
    2941.6336640213, 
    2718.91876032998, 
    2458.4890950268, 
    2326.39150999358, 
    1966.73139334906, 
    1882.46208246792, 
    1929.83996584002, 
    2071.27248705225, 
    1992.96095692882, 
    1729.78607224343, 
    1460.15786482461, 
    1293.93248942924, 
    1002.93947091681, 
    1101.71072201855, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    705.815881554449, 
    1280.47402830689, 
    1356.44093698884, 
    1398.61536541226, 
    1551.10838206687, 
    1699.38218059021, 
    1877.43620214529, 
    2156.54059274467, 
    2159.65305223428, 
    2208.47238213749, 
    2484.24128455779, 
    2376.76762415448, 
    2452.13636797355, 
    2520.54163015856, 
    2654.52729558819, 
    2647.2940070604, 
    2676.10395948489, 
    2712.18671056644, 
    2694.34172307483, 
    2824.03823525858, 
    3073.29597882659, 
    3109.38572266284, 
    3087.62761332142, 
    2993.08221813767, 
    3024.99009878861, 
    3061.06974626804, 
    3071.19122492722, 
    3062.79279038035, 
    2928.82844974626, 
    2710.74264508152, 
    2578.71856778211, 
    1891.99512387536, 
    2084.92961396778, 
    2154.77595364191, 
    2199.37708536626, 
    2229.32001731255, 
    1979.76314483143, 
    1874.21811542894, 
    1461.07034063063, 
    1013.3848108101, 
    760.115244378693, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    860.433289102615, 
    926.919156979619, 
    1156.44038810966, 
    1513.1839263256, 
    1599.08433148556, 
    1655.7181019003, 
    1911.80756535475, 
    2156.20961409112, 
    2212.91738160388, 
    2287.18595852627, 
    2337.64699483604, 
    2363.31183276097, 
    2582.34057959449, 
    2635.41094782779, 
    2656.29154062207, 
    2651.77663753181, 
    2660.27772386543, 
    2728.66792128572, 
    2827.29578688404, 
    2857.75619032425, 
    2975.76926251299, 
    3032.93980423934, 
    2995.5234596956, 
    3032.90651865624, 
    3085.86897090425, 
    3130.33488407758, 
    3194.49920930745, 
    3207.68038985466, 
    3041.10041494038, 
    2954.22772661489, 
    2693.34164275222, 
    2377.9294316204, 
    2374.25912464837, 
    2499.43204887163, 
    2473.5337632399, 
    2329.2342347008, 
    2011.64761229827, 
    1826.83408164901, 
    1496.49087953993, 
    1208.54294164573, 
    817.244186022817, 
    575.355392766152, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    787.652253490182, 
    991.559597834682, 
    1152.13735731784, 
    1364.85852264461, 
    1476.06714327115, 
    1451.2694311515, 
    1564.15081763172, 
    1850.86123159707, 
    2008.95865886639, 
    2132.17027990842, 
    2405.07124375232, 
    2466.32183982798, 
    2423.03918108799, 
    2578.84571758458, 
    2664.76363486543, 
    2652.36241937909, 
    2682.16524759646, 
    2665.47951178347, 
    2832.5265002374, 
    2939.95312244799, 
    2932.07698218348, 
    3041.37418959491, 
    3018.57197528027, 
    3003.75250988332, 
    3049.99118421886, 
    3102.92799160236, 
    3110.82732612087, 
    3066.83446804423, 
    3057.75541215554, 
    3034.00066651239, 
    2991.07887945701, 
    2895.11213049931, 
    2749.98800651536, 
    2657.48227873703, 
    2652.65663788299, 
    2519.09193871228, 
    2360.69310598777, 
    1973.96307423014, 
    1699.5520219145, 
    1894.90837449535, 
    1579.85833537298, 
    1081.99684031905, 
    491.518998346181, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1010.46756837054, 
    1185.8531365651, 
    1273.27715647828, 
    1547.20513043916, 
    1461.62480341715, 
    1504.97373300991, 
    1721.85181412918, 
    1929.16203307368, 
    2146.05045844658, 
    2204.051994343, 
    2189.8167210267, 
    2361.61233986136, 
    2493.95253805737, 
    2504.00274476191, 
    2633.0812443268, 
    2662.64214604814, 
    2700.43033499992, 
    2823.05235716393, 
    2874.68804217602, 
    2910.47838416339, 
    3020.3466293377, 
    3051.6885389016, 
    3047.23008624497, 
    3082.35527834545, 
    3145.03691975703, 
    3130.46445338971, 
    3014.03481350858, 
    2997.56480978095, 
    3015.40277003175, 
    3057.09743717091, 
    2962.4445037966, 
    2838.85297989128, 
    2726.36524703261, 
    2639.10503342318, 
    2506.44089393235, 
    2297.94956171073, 
    2069.6953124313, 
    1651.80056829564, 
    1387.5805822332, 
    1472.56956781723, 
    1095.74748181477, 
    844.390416750522, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    859.037831700638, 
    1191.54939721284, 
    1212.31193243353, 
    1347.95322739959, 
    1454.9383615632, 
    1509.66541078347, 
    1650.93023106697, 
    1918.2738499276, 
    2181.84814442332, 
    2210.66290468329, 
    2221.7813634193, 
    2454.1358705457, 
    2611.51961811489, 
    2579.61154130676, 
    2611.52616785027, 
    2687.57772003224, 
    2763.75309241053, 
    2781.23716052744, 
    2822.95051843694, 
    2868.65229344387, 
    2925.46599147951, 
    3048.82920800814, 
    3094.85732075386, 
    3129.48468658361, 
    3166.43563674419, 
    3171.8713431545, 
    3181.57673912319, 
    3017.60322875523, 
    3030.55372893377, 
    2957.38150123716, 
    2914.19221226314, 
    2834.20210283451, 
    2745.87799755613, 
    2627.88280990576, 
    2514.7808054506, 
    2345.38106432177, 
    2019.5905199342, 
    1674.67453047131, 
    1373.73187672065, 
    1420.55014655578, 
    1234.77133300299, 
    1430.29787020874, 
    1084.0854802214, 
    927.388263511814, 
    1580.53480216718, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    859.156334869042, 
    1099.82160903586, 
    1396.41943161818, 
    1514.20099450758, 
    1502.08053034084, 
    1760.01604173063, 
    1951.11636274229, 
    2116.07681488876, 
    2206.42534735513, 
    2299.65749529634, 
    2571.64023029651, 
    2756.49436067854, 
    2713.68877318958, 
    2677.37686514912, 
    2753.60120217509, 
    2810.86017048777, 
    2916.74575654397, 
    2984.04641718953, 
    2885.47036209929, 
    2904.74125888827, 
    3117.24690230224, 
    3136.4693074357, 
    3155.61476114238, 
    3162.30638025956, 
    3181.14317123005, 
    3170.13095962036, 
    3115.73722720127, 
    3124.93053363694, 
    3083.38980773875, 
    2982.28542572314, 
    2942.56514002044, 
    2774.42393708881, 
    2646.12427506721, 
    2424.77690019723, 
    2239.63344525677, 
    2028.86658758426, 
    1801.31226441421, 
    1477.09130616895, 
    1180.6852050774, 
    1290.4168105949, 
    1017.20673697308, 
    1827.08501040168, 
    587.923696398954, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1223.94850794876, 
    1258.18162539679, 
    1219.62589161034, 
    1309.54044338797, 
    1570.29519961466, 
    1660.93735571507, 
    1786.63619461201, 
    1928.89518871919, 
    2126.53646136627, 
    2220.8429538079, 
    2309.16407927628, 
    2601.07431903228, 
    2778.23396198124, 
    2701.80547961764, 
    2709.28322501239, 
    2761.73225172846, 
    2797.99018356035, 
    2943.81457350341, 
    3053.62852053893, 
    2963.59350263706, 
    3031.74629001717, 
    3123.24086722201, 
    3150.76331789418, 
    3158.72919959859, 
    3162.53418355409, 
    3118.07252953574, 
    3147.11430344344, 
    3134.08088457776, 
    3121.26796664685, 
    3136.81589135228, 
    2978.85455734234, 
    2880.64154152568, 
    2842.70218443076, 
    2694.14396316702, 
    2396.01128537213, 
    2251.24349445328, 
    2110.6749862173, 
    1935.97944961473, 
    1627.2885342293, 
    1350.73304394776, 
    1192.70979267084, 
    992.427451814946, 
    1348.10059549126, 
    2068.57261198104, 
    1304.13629241178, 
    1541.91912192344, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1224.37675931769, 
    1093.09944484562, 
    1269.78315179927, 
    1640.86105590611, 
    1638.71508575635, 
    1781.34621178048, 
    1953.36814564579, 
    2215.80129453108, 
    2309.43151473553, 
    2256.67349979669, 
    2409.26316428924, 
    2614.75760682362, 
    2684.47760626112, 
    2723.36767901865, 
    2790.59016569941, 
    2902.16059751529, 
    3017.16670799465, 
    3029.83164235482, 
    3071.92706037918, 
    3107.37465441583, 
    3082.42641071415, 
    3086.13299086218, 
    3150.14325320357, 
    3101.12380536437, 
    3123.4351562284, 
    3077.41799881276, 
    3023.70566396402, 
    3112.98688869768, 
    3084.3244489138, 
    2931.23219318233, 
    2878.25046331514, 
    2808.59955288105, 
    2684.55706528474, 
    2625.23817963211, 
    2417.32716528461, 
    2245.98921168986, 
    2005.01855200746, 
    1753.62762524574, 
    1811.3343397905, 
    887.218731686432, 
    1281.60571384927, 
    700.050673252336, 
    938.190634376819, 
    1706.87014070522, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1453.66870780441, 
    1085.94537455139, 
    1214.40367978384, 
    1559.80942088505, 
    1649.96520331846, 
    1920.7140527706, 
    2058.29586840885, 
    2346.96444387648, 
    2198.68665545228, 
    2173.91638123041, 
    2378.57982865988, 
    2556.11663093191, 
    2673.2568398224, 
    2774.77582174698, 
    2793.7781624155, 
    2908.56629695302, 
    2937.35136939902, 
    2964.23468487569, 
    3031.89937032491, 
    3013.53227067023, 
    2941.40762080123, 
    3007.9377004175, 
    3068.95727329762, 
    3081.13336807673, 
    3113.69200368765, 
    3108.40498956869, 
    3021.37329111541, 
    3075.44755919492, 
    3008.84012253793, 
    2918.70589389018, 
    2983.2859670757, 
    2831.39343471604, 
    2590.93403474898, 
    2559.5567195421, 
    2456.61900401185, 
    2306.77477251813, 
    1990.20167508583, 
    1473.29158810311, 
    1433.75812433128, 
    1346.80382002351, 
    1981.37402280321, 
    1091.03718514966, 
    1320.66570032443, 
    1182.87132405668, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    510.080579414127, 
    844.50256259262, 
    1005.97808799039, 
    979.051167878176, 
    1475.83976938477, 
    1461.65591518564, 
    1673.49562196741, 
    1866.31833684792, 
    2017.2092273751, 
    2278.37959790848, 
    2231.14225478252, 
    2271.88387361566, 
    2382.18586073585, 
    2521.72619622463, 
    2642.54538309337, 
    2736.23403552617, 
    2766.25462907472, 
    2871.21050844663, 
    2904.35099447142, 
    2957.75317461527, 
    3006.02528113155, 
    3074.86093951353, 
    3085.35898980686, 
    3032.53467616377, 
    3089.24102789929, 
    3145.95296495137, 
    3124.11785941118, 
    3108.38402180646, 
    3079.30317668354, 
    3006.34249752687, 
    2984.87032688507, 
    2931.76969748518, 
    2821.45116044666, 
    2776.76211132227, 
    2603.32695547076, 
    2508.1589408047, 
    2431.66699592046, 
    2339.6446563653, 
    2015.21932536737, 
    1398.18299515488, 
    1160.92649873472, 
    927.684708660972, 
    1002.96047971852, 
    1036.68433365646, 
    903.110278602388, 
    965.772626661171, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    863.532443121153, 
    869.337359404157, 
    1214.724014411, 
    1492.16739021439, 
    1637.50417504324, 
    1782.00656029545, 
    1996.56615463103, 
    1928.12066321935, 
    2041.69489989381, 
    2278.06215166803, 
    2458.27450730563, 
    2479.68378510237, 
    2623.52896942177, 
    2715.92510418131, 
    2796.77310262873, 
    2852.86032771573, 
    2947.25959502727, 
    3026.79083597945, 
    3044.44421521019, 
    3123.99251875609, 
    3151.50491279794, 
    3114.21984733732, 
    3186.87792826449, 
    3281.85999304944, 
    3202.040127748, 
    3097.21695737736, 
    3126.22810858511, 
    3056.29465234186, 
    3006.6003496977, 
    2952.35352748916, 
    2794.48530764367, 
    2656.57290662715, 
    2654.63345036754, 
    2563.98758678032, 
    2425.64957649184, 
    2355.44557083582, 
    2163.07997335125, 
    1711.88901809598, 
    1070.67904958466, 
    887.727004815499, 
    991.930789435443, 
    1004.73041283892, 
    953.379570150075, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    917.462256557567, 
    1253.04501057811, 
    792.658455315077, 
    1165.59741837664, 
    1327.4823397507, 
    1559.91377699019, 
    1582.45420315864, 
    1799.38146121656, 
    1979.84557247123, 
    2011.35352534892, 
    2065.50900810405, 
    2267.89690598393, 
    2379.44678350557, 
    2468.55034658818, 
    2598.63389815957, 
    2771.18604633038, 
    2860.63645033357, 
    2925.93048230926, 
    2942.22584333304, 
    3033.70466115848, 
    3137.25795841269, 
    3160.4774033207, 
    3187.74537345804, 
    3286.10917804702, 
    3344.02178228476, 
    3369.55632393716, 
    3204.04634197684, 
    3270.664141768, 
    3222.31757616559, 
    3089.00006013079, 
    3124.53994576556, 
    2994.87860685624, 
    2929.85264683609, 
    2782.46864439927, 
    2701.45554899259, 
    2588.63603023755, 
    2540.97316637919, 
    2396.54019567681, 
    2046.93208601223, 
    1786.82928921946, 
    1862.04413564227, 
    976.858502691464, 
    1293.30287199949, 
    568.035233827688, 
    735.145546364845, 
    0, 
    623.184348865827, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    778.359072420551, 
    1035.7482548919, 
    833.193083042089, 
    1140.64267115725, 
    1535.11499711021, 
    1356.36642096521, 
    1638.6090277157, 
    1920.93613325331, 
    2086.05430902196, 
    2152.38127025147, 
    2351.39882328795, 
    2520.14553451792, 
    2561.24747890955, 
    2647.58575669962, 
    2830.5202448468, 
    2927.93026938936, 
    2991.93566430039, 
    3062.57186211803, 
    3127.29950170805, 
    3194.49441228891, 
    3210.31724297245, 
    3242.32184320852, 
    3338.41897876643, 
    3373.18211277794, 
    3323.27939625862, 
    3231.54247558543, 
    3092.11755904091, 
    3053.09630189306, 
    2835.58377382007, 
    3000.61820933234, 
    2968.97725310885, 
    3029.45698251408, 
    2864.97542079724, 
    2792.71838769493, 
    2595.45682716055, 
    2358.83511093284, 
    2512.66076755686, 
    1914.63635678923, 
    1518.81417233899, 
    1406.9944272188, 
    1313.59846196683, 
    769.93881431295, 
    881.667404781102, 
    1240.13831813279, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    560.685172429394, 
    1074.35964442371, 
    1867.07090572274, 
    1833.36064965142, 
    1565.20874375918, 
    1645.08191977116, 
    2012.83848998527, 
    2266.89714508292, 
    2278.57118065854, 
    2404.684569706, 
    2510.6263193852, 
    2664.00551712029, 
    2793.61531204234, 
    2926.30792696148, 
    3023.92106341826, 
    3068.9083816918, 
    3122.74446107889, 
    3202.62323249418, 
    3253.54879127075, 
    3271.96794748409, 
    3256.58109730576, 
    3278.66632811601, 
    3292.73558989254, 
    3348.67875730912, 
    3316.23870885872, 
    3145.98263201903, 
    2776.45942573421, 
    3004.67763242245, 
    2863.16262716898, 
    2846.89145841456, 
    2916.84908530726, 
    2917.05811811697, 
    2848.05506398863, 
    2724.80244468942, 
    2294.0517317839, 
    2002.90904104757, 
    1761.53492297931, 
    1120.99119610366, 
    1179.20911560977, 
    968.205585017788, 
    1494.40367285638, 
    845.043548666602, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    561.535710463896, 
    1843.79724277119, 
    1586.98660837191, 
    1496.07142611015, 
    1680.37425946659, 
    1843.3319639877, 
    2104.61508304198, 
    2323.74795108018, 
    2342.78243536297, 
    2487.25131521845, 
    2557.46227921829, 
    2736.61410744685, 
    2892.21813410562, 
    3010.73732980961, 
    3098.50574194024, 
    3105.66195869934, 
    3168.132364813, 
    3235.46466989747, 
    3255.20521859632, 
    3245.05406208194, 
    3256.24564407863, 
    3220.00383697964, 
    3186.62931213992, 
    3124.99179953982, 
    3130.84826000324, 
    2952.32150574812, 
    2772.82689663484, 
    2730.43810129463, 
    2817.87874134683, 
    2710.02584907963, 
    2773.34379290133, 
    2800.30353925643, 
    2833.80685535449, 
    2810.45059859335, 
    2282.59565004058, 
    1826.68858017221, 
    1812.74274443281, 
    1351.48721584144, 
    1547.94324210786, 
    1066.56917559424, 
    1508.34982382989, 
    1784.79233088328, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    928.661915199837, 
    963.357251542481, 
    1048.71141453187, 
    1386.4377661331, 
    1620.38984643894, 
    1933.96599700007, 
    2074.57994632734, 
    2186.13906756107, 
    2299.55812506582, 
    2459.87555401668, 
    2601.89805674321, 
    2748.20770933913, 
    2883.53736570981, 
    3012.69406938975, 
    3095.1471937958, 
    3135.91863602314, 
    3209.71502846781, 
    3227.30511955546, 
    3234.08006288756, 
    3212.79114288552, 
    3216.42664849262, 
    3199.15685324337, 
    3113.62085741716, 
    3084.90745292798, 
    3129.11566041035, 
    2980.9823952211, 
    2778.97136474012, 
    2585.60699991104, 
    2593.17034975459, 
    2615.69971443012, 
    2695.67635567204, 
    2518.78724192019, 
    2644.45726718028, 
    2732.59915904673, 
    2615.67385190608, 
    2005.14430069548, 
    1722.19530306256, 
    1306.93026766626, 
    1337.16244566359, 
    998.088925170709, 
    1004.95870177713, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    443.957651509719, 
    1042.66831333721, 
    1246.13227264881, 
    1535.35395497226, 
    1822.14395193175, 
    1841.89809851696, 
    1963.62019101651, 
    2047.93869517265, 
    2181.58575377228, 
    2487.95789449171, 
    2675.63741370325, 
    2752.23352682101, 
    2844.48296319616, 
    2943.34963422439, 
    3065.89081231115, 
    3233.32637580981, 
    3137.46241595304, 
    3146.45822718149, 
    3198.6875642102, 
    3077.6132687128, 
    3156.43476379242, 
    3138.52106248875, 
    3087.49625163158, 
    3099.14860221623, 
    3101.26943249001, 
    3038.07036832327, 
    2870.37007041973, 
    2716.54449687007, 
    2537.77548844418, 
    2639.25084125706, 
    2738.88897183059, 
    2663.97546642879, 
    2681.87779412926, 
    2648.30055184068, 
    2624.80056137775, 
    2446.44229878224, 
    1936.87319242652, 
    1565.95187705647, 
    1593.02613914432, 
    1259.65053036594, 
    753.683659332421, 
    671.528665688685, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    626.541329803487, 
    562.712095569241, 
    983.781550821181, 
    1135.46558422554, 
    1342.14565082916, 
    1754.20771326957, 
    1799.08021589626, 
    1822.39193427929, 
    1859.02251465952, 
    1963.67665909177, 
    2214.78490949224, 
    2453.88832928061, 
    2618.37124562289, 
    2748.32197597503, 
    2873.59290228528, 
    2959.50714847628, 
    3091.52878942352, 
    3035.33799496064, 
    3175.41308660007, 
    3242.88914961368, 
    3146.58072742131, 
    3117.92366056988, 
    3149.51702268482, 
    3180.34725541042, 
    3162.24898615907, 
    3112.63421338492, 
    3069.79430435426, 
    3031.0774310681, 
    2960.18033373038, 
    2822.08660918501, 
    2479.04681665911, 
    2413.10795042314, 
    2688.81656769425, 
    2648.65519779071, 
    2434.41045779832, 
    2461.32382826926, 
    2234.26746508528, 
    2082.34922489291, 
    1786.37821018563, 
    1478.50745751014, 
    1209.52723873219, 
    1265.8046685589, 
    1174.60003944001, 
    1069.715561902, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    558.194521089731, 
    907.155754072977, 
    1222.18539225669, 
    1447.329368952, 
    1710.34730164235, 
    1652.35781154749, 
    1775.09029140625, 
    1826.93681840642, 
    1852.78453287832, 
    2232.90573816856, 
    2460.22520987549, 
    2626.87324828105, 
    2749.27550563974, 
    2910.19435471178, 
    3080.5626178281, 
    3165.67170233494, 
    3107.06643360826, 
    3190.33476332648, 
    3236.59479970819, 
    3135.26981670956, 
    3091.51731000977, 
    3077.34723999007, 
    3187.42004188657, 
    3142.12355967024, 
    3163.35046974786, 
    3223.22263470266, 
    3092.3484617345, 
    3000.92691623251, 
    2835.21856818573, 
    2437.00468353129, 
    2137.6387240505, 
    2203.03067467175, 
    2406.00242829367, 
    2294.21838410104, 
    2239.74494252103, 
    2261.19506059524, 
    1995.96398419403, 
    1866.17122356571, 
    1571.33835070377, 
    1269.06965141428, 
    974.020737256273, 
    1323.87080111375, 
    896.178992533862, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    693.817830618458, 
    706.950454252287, 
    806.37703442659, 
    962.384332933729, 
    1224.34754396717, 
    1309.64773500415, 
    1531.49925305127, 
    1721.56070097517, 
    1671.99899010397, 
    1791.61600386172, 
    1904.57165236745, 
    2067.14503699304, 
    2339.02031825583, 
    2460.68326798666, 
    2559.72349471998, 
    2731.77972336333, 
    2879.62754044477, 
    3042.05094271118, 
    3186.63085209984, 
    3141.11578120801, 
    3211.54454821536, 
    3168.45598234534, 
    3146.41039259128, 
    3109.47297588168, 
    3074.76416958802, 
    3092.88899228681, 
    3108.60061457735, 
    3142.386172051, 
    3177.85870219628, 
    3160.73928930392, 
    3037.52934072119, 
    2715.47779281378, 
    2456.03840314196, 
    2300.95605058006, 
    2399.61984183862, 
    2434.93342100685, 
    2158.39061619765, 
    2113.66956372501, 
    2167.14424957176, 
    1656.40799439241, 
    1505.30007517229, 
    1766.80659721062, 
    903.528674472162, 
    491.021686924717, 
    0, 
    1313.20177133654, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    690.299686956574, 
    1031.36917649373, 
    1088.89170208798, 
    1203.98581205431, 
    1269.84740187719, 
    1401.19468362397, 
    1520.56351241581, 
    1580.45917319583, 
    1565.46667998642, 
    1708.53781867055, 
    1889.74550783206, 
    2027.73363607939, 
    2240.79196283044, 
    2456.82734234127, 
    2520.74792336119, 
    2608.88020599415, 
    2703.33999641712, 
    2819.61626942528, 
    2987.57718251476, 
    3157.7316904421, 
    3179.38166252658, 
    3141.06501445077, 
    3158.12428722298, 
    3173.48085596594, 
    3249.38901456556, 
    3185.12727522224, 
    3159.38114042269, 
    3115.19394007027, 
    3139.4738876094, 
    3127.13447052589, 
    3168.37780244692, 
    2978.47051278434, 
    2519.28949691716, 
    2620.42996377875, 
    2492.56936767845, 
    2587.56261836053, 
    2266.28967329263, 
    1980.57561106169, 
    2059.52843531467, 
    2230.27263713341, 
    1482.50795329399, 
    1641.73121345754, 
    1096.3777451619, 
    835.478333511695, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    556.21661134006, 
    794.885278483855, 
    0, 
    1354.15897725823, 
    1215.27036638714, 
    1279.3131569444, 
    1520.36390890193, 
    1612.80526505912, 
    1661.55442717106, 
    1655.87787878009, 
    1868.43831964229, 
    1994.06351014287, 
    2093.06820579392, 
    2286.82147074673, 
    2427.53038601418, 
    2480.19417737966, 
    2574.86634964704, 
    2669.57580498823, 
    2853.93842827438, 
    3002.13619949972, 
    3142.54546219838, 
    3249.51888125554, 
    3153.78933213948, 
    3167.34585714505, 
    3191.28256024392, 
    3148.61066785206, 
    3195.65003254129, 
    3224.3045449017, 
    3268.40474646885, 
    3219.48737608552, 
    3219.42581416306, 
    3104.15117192311, 
    2873.64692513496, 
    2747.31176327236, 
    2853.09652602598, 
    2595.39229587252, 
    2330.79211703697, 
    2081.52523852203, 
    1926.04833962891, 
    1911.91258336899, 
    1838.07255944108, 
    1440.05318488861, 
    1345.82214371979, 
    690.243644867299, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    970.987707001602, 
    963.650419850129, 
    994.981555388217, 
    1156.06364277901, 
    1311.2636721261, 
    1477.3788649852, 
    1622.66937965798, 
    1747.26220701933, 
    1699.94631879219, 
    1860.97460517822, 
    2001.69127373897, 
    2107.07240240994, 
    2255.23762014954, 
    2464.63478906818, 
    2568.98032721113, 
    2648.71564057396, 
    2754.54774890689, 
    2864.21532387287, 
    2948.56126190248, 
    3156.63321381212, 
    3363.50127575825, 
    3177.58101444124, 
    3163.66590477999, 
    3229.66843771177, 
    3272.65318736983, 
    3243.27697573287, 
    3255.86136790835, 
    3320.67538196374, 
    3291.42373135322, 
    3083.87946004568, 
    3029.16036482555, 
    3119.29871927525, 
    2690.13041158645, 
    2597.05295992623, 
    2544.36539453167, 
    2403.8892827577, 
    2049.58905545608, 
    2076.30278154853, 
    1755.98882040548, 
    1933.61476719081, 
    1334.21016118098, 
    1023.80049725791, 
    832.114285070855, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    981.222077729342, 
    1047.33193656888, 
    1086.30662102062, 
    1205.76675402047, 
    1424.03370852712, 
    1484.09778407302, 
    1568.22167470768, 
    1619.2413928836, 
    1703.69381050693, 
    1853.64725157296, 
    1989.67595027063, 
    2133.57966447694, 
    2225.90896866772, 
    2397.31758839723, 
    2560.62001080075, 
    2705.83439886182, 
    2755.10653334972, 
    2850.00773654598, 
    2943.2110185841, 
    3088.90761960295, 
    3312.07921255958, 
    3192.20149990563, 
    3208.58737205032, 
    3282.13588042152, 
    3313.86756991869, 
    3344.12047333401, 
    3320.72017696503, 
    3323.71321864536, 
    3304.3302862929, 
    3002.15083776113, 
    2971.95193455358, 
    2991.31378233865, 
    2823.66512933663, 
    2468.03171584535, 
    2588.8954975777, 
    2650.16152174703, 
    2426.23931856806, 
    1991.21338793579, 
    2003.30585891641, 
    1884.07979636185, 
    1386.5488393971, 
    1167.32527685031, 
    789.257360405196, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    950.765787383883, 
    1100.54774866811, 
    1133.14769216996, 
    1315.1476816163, 
    1485.23322637578, 
    1436.32521588428, 
    1538.50191502947, 
    1640.37731992084, 
    1678.6162723074, 
    1838.83303818146, 
    1968.5062323456, 
    2123.81773256706, 
    2200.59601651104, 
    2353.51022300229, 
    2510.16378232784, 
    2618.34182790894, 
    2738.59606670547, 
    2864.27971758189, 
    2920.3054842482, 
    3065.67040700858, 
    3212.60404595432, 
    3225.54908708513, 
    3238.55705126864, 
    3314.51084126761, 
    3330.68889231531, 
    3352.88752998838, 
    3388.32935106121, 
    3231.79966565855, 
    3248.71108775285, 
    3130.73155763945, 
    3134.7295424756, 
    3230.86786120774, 
    2837.13431280256, 
    2417.99527971312, 
    2689.36680744497, 
    2882.6052012779, 
    2653.65689632772, 
    2178.19502825456, 
    2337.34141692611, 
    2095.69221967405, 
    1602.35400352816, 
    1412.10425586241, 
    700.544265798805, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1000.52815000693, 
    1053.84529616061, 
    1393.52904607351, 
    1654.87089809246, 
    1485.41568648306, 
    1524.68089491838, 
    1573.72468337811, 
    1665.72702439428, 
    1926.98885184059, 
    1972.97189332014, 
    2110.35421809884, 
    2222.83531382826, 
    2414.8142284162, 
    2503.52338680785, 
    2577.61843250812, 
    2728.66617920079, 
    2809.298532839, 
    2909.75023392144, 
    3032.38693112655, 
    3100.70261430325, 
    3141.14478805432, 
    3236.92892572063, 
    3295.2908041922, 
    3329.78709512643, 
    3327.57264814017, 
    3293.87030760535, 
    3037.22779107404, 
    3117.26698523423, 
    3268.96640440484, 
    3233.7456492479, 
    3130.22476444688, 
    2898.34862702654, 
    2488.86465950764, 
    2988.39488846441, 
    2627.64055528823, 
    2033.3845991579, 
    1970.80639732424, 
    2302.82885418665, 
    2275.49401197948, 
    1591.2487675698, 
    1154.63036028815, 
    914.695730137693, 
    739.290480371364, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    933.217284258756, 
    1018.92800953574, 
    1027.35511695593, 
    1323.02566018321, 
    1583.86915840139, 
    1589.43795074726, 
    1604.57514662597, 
    1627.07925755238, 
    1690.71976184107, 
    1946.01307976237, 
    2042.76140001913, 
    2130.36110745886, 
    2240.48287034048, 
    2412.07210691095, 
    2546.8613392519, 
    2656.3808043869, 
    2783.38771034315, 
    2842.0695223452, 
    2914.31533957516, 
    2996.56037609084, 
    3067.46096848942, 
    3154.5893339382, 
    3260.64837854658, 
    3300.05795926291, 
    3303.00287515612, 
    3283.5570363649, 
    3243.59782619409, 
    3150.21395235596, 
    3098.37249870873, 
    3184.31328643767, 
    3216.38713045286, 
    3179.81742870946, 
    2945.62718942794, 
    2866.35054711498, 
    3015.21995625953, 
    2588.34443890858, 
    2109.18568704126, 
    2019.61914390857, 
    2439.91665465383, 
    2189.34921594255, 
    1581.72713503592, 
    1332.31127272666, 
    1157.29258758291, 
    865.678224742982, 
    750.336112262388, 
    882.431727454513, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    776.114189491349, 
    1077.15565730559, 
    1029.50483146857, 
    1338.30906265108, 
    1552.65059090296, 
    1637.87538317044, 
    1672.40327873095, 
    1655.54317661177, 
    1772.86030153972, 
    1881.5193924087, 
    1966.64016078662, 
    2148.28442002379, 
    2307.64831949894, 
    2418.8057077693, 
    2556.58539417412, 
    2596.13217764728, 
    2648.73358969464, 
    2833.98699580597, 
    2922.53682300254, 
    2981.43450626499, 
    3063.18883695866, 
    3171.97806954426, 
    3223.5019541407, 
    3245.87758333579, 
    3259.04731169717, 
    3205.92164599963, 
    3189.48628734885, 
    3215.04626928103, 
    3182.92888261784, 
    3171.99181456782, 
    3102.82394773233, 
    3044.94231253398, 
    2840.59114638411, 
    2782.50784343795, 
    2980.35167072866, 
    2588.96727664699, 
    2243.86157756433, 
    2287.23019819577, 
    2307.22820984303, 
    1907.99925903729, 
    1758.59197294532, 
    1487.51956316456, 
    1346.23932291113, 
    1297.5490671897, 
    995.043746816778, 
    913.668073141133, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    932.334322091572, 
    1050.32562828208, 
    1506.9452306057, 
    1542.22513749391, 
    1655.37629616092, 
    1661.92754812944, 
    1632.83892154245, 
    1685.13345203901, 
    1775.70903808886, 
    1940.04632932857, 
    2165.80689140609, 
    2322.75251698342, 
    2496.68808561266, 
    2545.75485378233, 
    2508.25254763834, 
    2553.57349833918, 
    2743.60958951583, 
    2885.21776486295, 
    2946.77906717148, 
    3039.41424773152, 
    3189.58756812517, 
    3215.54639302276, 
    3208.8229432396, 
    3189.52316451326, 
    3180.54239072455, 
    3171.92099305535, 
    3155.35766319969, 
    3136.59096113421, 
    3030.87812836702, 
    3105.77003797784, 
    3080.14529300432, 
    2984.40773181209, 
    2776.70631567513, 
    2702.78673771268, 
    2527.93683701388, 
    2249.80948767741, 
    2547.0912526998, 
    2336.77251157179, 
    2075.59581732301, 
    1752.63805660734, 
    1482.09991702656, 
    1292.93775565639, 
    1224.68583889528, 
    1149.57842782406, 
    919.65316886397, 
    836.086596209797, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    961.890367385508, 
    1174.23407804214, 
    1274.79598272904, 
    1348.49945000969, 
    1620.55849261097, 
    1565.73263680351, 
    1703.70236285794, 
    1773.74545223715, 
    1715.97002049941, 
    1849.95532375782, 
    2056.28199566075, 
    2251.52822997403, 
    2404.53309169214, 
    2416.59744924012, 
    2492.81247485031, 
    2594.48345971266, 
    2743.82219315929, 
    2848.00607514736, 
    2938.19511374689, 
    3044.91759042677, 
    3248.12341681299, 
    3188.69927223366, 
    3194.93272416112, 
    3123.33497203685, 
    3122.03547083416, 
    3115.46131520517, 
    3103.63138004109, 
    3201.73483884981, 
    3086.8080263794, 
    3100.90801504241, 
    3096.53112845203, 
    2879.46842643035, 
    2585.63122757658, 
    2552.0042603625, 
    2612.24161128434, 
    2591.1757458112, 
    2602.55561207226, 
    2435.91524011292, 
    2100.28150306782, 
    1921.3450548308, 
    1762.81758274343, 
    1471.35936274966, 
    1274.33038137823, 
    1639.06709796729, 
    1250.62393080543, 
    710.292792272106, 
    576.884354181355, 
    462.164874383782, 
    968.291038132256, 
    947.972227313993, 
    511.13487742568, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    891.301341402766, 
    1030.8971023948, 
    1226.45892360817, 
    1265.88926889774, 
    1336.03198624033, 
    1525.05367214133, 
    1515.52680225507, 
    1668.55225072324, 
    1637.98886487036, 
    1615.62639250165, 
    1786.06566331643, 
    2021.79132122915, 
    2231.62212966932, 
    2366.59585551591, 
    2369.17080442157, 
    2510.42356794883, 
    2684.69270775488, 
    2764.71188623132, 
    2828.55576730632, 
    2925.09162282878, 
    3060.4018216087, 
    3248.70598901157, 
    3176.64685116487, 
    3187.60234835807, 
    3148.86649491268, 
    3145.71168682241, 
    3146.80789560519, 
    3057.80198151324, 
    3049.22228980071, 
    3053.03573678586, 
    3119.76570984845, 
    2979.16624684321, 
    2658.10331488712, 
    2569.56100407061, 
    2453.01962011846, 
    2530.20365398327, 
    2605.60542802409, 
    2564.837431152, 
    2498.2143903234, 
    2358.48427823429, 
    2275.66680281199, 
    1894.53143892611, 
    1561.90099728738, 
    1616.07396674255, 
    1458.19338644878, 
    1376.07625502418, 
    1124.81451121174, 
    1024.87200241448, 
    1224.03811047505, 
    1226.07811084381, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1069.08664851413, 
    1190.49040819932, 
    1326.45156751976, 
    1410.92202305585, 
    1582.6286642675, 
    1424.86151436145, 
    1467.45571441434, 
    1562.04989030703, 
    1649.46835732687, 
    1751.70498571953, 
    1987.45190950605, 
    2220.18524331783, 
    2329.33414785972, 
    2332.4898411549, 
    2553.92712650905, 
    2752.38838715673, 
    2744.22540026696, 
    2828.74114140902, 
    2925.9751906555, 
    3102.43025296191, 
    3152.60837107152, 
    3143.33506052514, 
    3160.98860252718, 
    3148.6092239896, 
    3109.90179633559, 
    3135.39161345846, 
    3116.30361222733, 
    3104.17174119648, 
    3195.67869097139, 
    3193.31181592509, 
    3045.37965792453, 
    2787.34669718457, 
    2584.72461849487, 
    2482.68220375503, 
    2402.57295350686, 
    2360.76556109755, 
    2313.99953247821, 
    2404.50325574979, 
    2377.39855419038, 
    2447.83225448654, 
    2148.64953592678, 
    1772.85260638204, 
    1729.02764231833, 
    1878.3352373936, 
    1679.91719446771, 
    1519.37997819201, 
    1141.06976531101, 
    1462.1290920368, 
    1112.12951692774, 
    491.361055742664, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    900.265082534727, 
    1118.48788633601, 
    1101.36567604628, 
    1345.3681465211, 
    1406.82892330754, 
    1456.95263910247, 
    1444.15592245277, 
    1561.94268030111, 
    1715.59371326356, 
    1790.11275879285, 
    1948.98920725359, 
    2029.91687461041, 
    2200.29724243882, 
    2286.10456586741, 
    2420.63306564956, 
    2660.93989380008, 
    2702.98712142373, 
    2758.45580554789, 
    2877.26963170734, 
    3024.03502151234, 
    3124.47208578571, 
    3124.52218661458, 
    3144.15471784464, 
    3141.39840867861, 
    3142.94335466099, 
    3142.56499278228, 
    3092.52732300472, 
    3191.78922623444, 
    3161.83559491591, 
    3140.22555549184, 
    3105.25605465904, 
    3070.85383954424, 
    2839.55984286107, 
    2716.69653830245, 
    2504.48922693627, 
    2287.65182152665, 
    2303.81556882481, 
    2335.59206808358, 
    2387.7958984042, 
    2208.03818705145, 
    2136.93548178428, 
    2022.33321134921, 
    1918.0918558898, 
    1837.96974275525, 
    1721.95357372869, 
    1575.58666590575, 
    1145.8947185748, 
    1139.1217076918, 
    1164.33352733256, 
    818.409000092103, 
    492.044519352939, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1015.26163874829, 
    1243.1487074315, 
    1423.94430891866, 
    1385.95892038968, 
    1363.37954985966, 
    1419.73348316989, 
    1594.30709549619, 
    1796.10301327541, 
    1978.85603586653, 
    2097.04133358051, 
    2116.4551275694, 
    2153.57031266761, 
    2320.67246712717, 
    2462.11703675889, 
    2686.37378697772, 
    2754.74026705094, 
    2788.7626130737, 
    2905.87771939769, 
    3059.35525621071, 
    3101.84276544885, 
    3129.8034802407, 
    3146.1246675904, 
    3143.2458690137, 
    3131.3923439532, 
    3099.03202864974, 
    3040.68629816739, 
    3071.59030137575, 
    3016.58641803105, 
    3009.75879958383, 
    3016.43551995446, 
    2963.86154791751, 
    2778.28128731904, 
    2683.34513101532, 
    2489.8269576384, 
    2286.76784316197, 
    2423.51088511546, 
    2337.10640180874, 
    2454.96443574108, 
    2235.79959918208, 
    2010.08061105559, 
    1996.88469188921, 
    1846.9594315336, 
    1754.74874717914, 
    1761.95492107794, 
    1746.02320828869, 
    1707.83747707859, 
    1399.26358669339, 
    1137.85824367194, 
    889.338913973714, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1070.09397800727, 
    1366.6806614523, 
    1341.49344091951, 
    1340.21203738842, 
    1385.20574940672, 
    1368.56036576708, 
    1557.29021557058, 
    1795.70828043705, 
    1951.84707939389, 
    1982.75157156038, 
    2118.47865548248, 
    2207.48273354627, 
    2160.04881015047, 
    2343.55791251623, 
    2483.11790789671, 
    2688.63186819555, 
    2853.58992231848, 
    2827.99420842054, 
    2908.6543227974, 
    3090.03286381311, 
    3064.86069539253, 
    3123.21779211479, 
    3121.38403238899, 
    3073.77250570215, 
    3074.5191632655, 
    3057.27795791525, 
    3006.95581535791, 
    3017.56750933536, 
    2892.12846248652, 
    2791.60524200251, 
    2811.38535188449, 
    2769.94325645479, 
    2665.47610429318, 
    2667.38021534111, 
    2489.27357311924, 
    2432.74487369865, 
    2531.78566015871, 
    2392.77173228159, 
    2379.25746112973, 
    2181.00231857522, 
    1865.83182127995, 
    1794.83151873627, 
    1596.92079072382, 
    1816.14833555776, 
    1457.71553258993, 
    1687.61356006601, 
    1778.11269948594, 
    1281.6628233646, 
    1069.09694622652, 
    556.402507920917, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1058.6031319665, 
    1142.99376978155, 
    1238.09751429449, 
    1312.56048463855, 
    1431.78024682096, 
    1419.23785319792, 
    1441.88396560575, 
    1535.7760630346, 
    1688.89455601325, 
    1917.78657389023, 
    2059.41146153906, 
    2032.33380028322, 
    2170.31834953954, 
    2317.47926470624, 
    2440.9509289641, 
    2621.44392552529, 
    2663.48114904617, 
    2779.19581020757, 
    2953.28171715926, 
    3092.52243593996, 
    3049.87075845084, 
    3122.15275063404, 
    3123.32807566223, 
    3096.64245765276, 
    3093.71059705521, 
    3050.38114693604, 
    2979.88770080137, 
    2939.09687068234, 
    2851.62387319074, 
    2769.26082273985, 
    2769.73799164193, 
    2756.35729676268, 
    2644.5291449299, 
    2703.60851601837, 
    2658.93445716255, 
    2612.15554053973, 
    2609.57024529766, 
    2437.04242794221, 
    2325.08497126086, 
    2132.82535272953, 
    2010.67622332279, 
    1887.53524396812, 
    1573.23158659558, 
    1774.87700629514, 
    1283.43450428842, 
    1185.3294689648, 
    1066.17919320331, 
    1349.60913548307, 
    995.494281936471, 
    416.127604499741, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    962.322332497751, 
    829.588944556798, 
    1120.29018958186, 
    1317.24119516365, 
    1380.09597480165, 
    1433.99263080764, 
    1625.28790082689, 
    1600.17073630896, 
    1754.80627615779, 
    1980.65570305266, 
    2159.41569186125, 
    2212.33968441895, 
    2304.6507347508, 
    2350.68945719176, 
    2434.73631528092, 
    2575.32908273817, 
    2679.5388086483, 
    2833.36847792246, 
    2960.7133529014, 
    3039.50579297311, 
    3063.74782837306, 
    3101.49401062567, 
    3083.41551102125, 
    3077.41965249824, 
    3094.87060138302, 
    3040.82695600312, 
    2966.85386928271, 
    2874.54488543524, 
    2787.26482902871, 
    2753.97538416827, 
    2775.23043654305, 
    2667.78654985517, 
    2708.20521577589, 
    2757.69651897979, 
    2803.6606907755, 
    2652.02645482248, 
    2543.40959974169, 
    2370.86641700648, 
    2379.78413800088, 
    2220.58597060934, 
    2006.86241186105, 
    1840.94057584632, 
    1735.14080479059, 
    1854.15561309493, 
    1032.60227739817, 
    594.543845651108, 
    838.304940931479, 
    1267.97227810368, 
    1508.53045056327, 
    735.365796902706, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1000.26421500956, 
    1257.13356055141, 
    1173.77262903856, 
    1297.07633416367, 
    1266.63677013375, 
    1423.25461686689, 
    1704.78068088668, 
    1811.80001111264, 
    1945.27162296799, 
    2005.95215892306, 
    2232.92069179683, 
    2401.08366387028, 
    2444.18276831857, 
    2500.42642629011, 
    2632.63122014437, 
    2814.38993310324, 
    2976.85963948495, 
    2946.36953645608, 
    3072.64171655253, 
    3123.02533633417, 
    3028.85814151659, 
    3053.14173351979, 
    3054.32733172731, 
    3069.1177365644, 
    3039.56977382712, 
    2939.2706310261, 
    2853.89705301307, 
    2786.41794284608, 
    2731.60494943596, 
    2661.07853495516, 
    2559.80043983, 
    2553.15149620432, 
    2684.13207581582, 
    2646.82844386229, 
    2406.70538276972, 
    2448.01668391968, 
    2442.28425989273, 
    2240.63805095664, 
    2189.86343734193, 
    2111.38082997549, 
    1947.89396242853, 
    1928.29242922188, 
    1327.67785104688, 
    831.968340796087, 
    0, 
    719.166992088221, 
    1485.40590846506, 
    1706.70566399903, 
    751.543598504944, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1109.93371973793, 
    1027.74386449292, 
    1225.93167119478, 
    1383.13858785016, 
    1388.80809200797, 
    1369.82891705805, 
    1427.62427982061, 
    1826.29077909799, 
    1837.42267800442, 
    1887.94576756676, 
    1971.52276101722, 
    2344.46265159591, 
    2432.61170794094, 
    2485.32127920246, 
    2559.03169217604, 
    2661.84536884401, 
    2696.13330499223, 
    2783.30271431657, 
    2921.85457070792, 
    2963.77785156339, 
    3028.96700919647, 
    3018.91441323623, 
    3045.77332107803, 
    3058.64406137453, 
    3052.45563617265, 
    2982.57587382291, 
    2853.93350203988, 
    2795.80164088718, 
    2714.16339355758, 
    2647.14799345699, 
    2618.74494579379, 
    2570.6740443066, 
    2504.78411171785, 
    2609.11823663971, 
    2696.44195334591, 
    2508.70573472343, 
    2415.01189714816, 
    2355.05497871028, 
    2155.51468089491, 
    2136.60491422112, 
    2003.63077230711, 
    1752.18836232858, 
    1438.67537359916, 
    740.421282869729, 
    716.500296488017, 
    0, 
    0, 
    998.083856562298, 
    1300.00211348342, 
    793.547996223469, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1074.69080864583, 
    992.884157225885, 
    1233.62477647889, 
    1353.56666833914, 
    1415.26669706433, 
    1521.12008075538, 
    1406.40256693071, 
    1548.52378265137, 
    1718.54353602279, 
    1845.27224119012, 
    1877.62735628429, 
    2160.53768226784, 
    2429.85014586049, 
    2498.49032915016, 
    2618.0165493968, 
    2673.42076306161, 
    2698.08415084758, 
    2761.81345371676, 
    2810.42929584451, 
    2896.88681215906, 
    2956.89457678697, 
    3073.87961064506, 
    3019.7718835027, 
    3061.63327995732, 
    3062.07399937683, 
    3071.08506039799, 
    2999.41775384875, 
    2841.67125654993, 
    2746.70352650095, 
    2696.08967524822, 
    2638.90743083589, 
    2607.32019174182, 
    2559.45199498786, 
    2520.5549900412, 
    2571.80430505203, 
    2518.3156549361, 
    2651.0806594068, 
    2519.57298067905, 
    2471.65614622191, 
    2288.84652525795, 
    2068.32560960807, 
    1912.80346432265, 
    1525.28875490727, 
    1511.28283296242, 
    1029.19930794597, 
    662.717912126677, 
    0, 
    0, 
    1036.11665405047, 
    1306.57355805547, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1121.52897057209, 
    1165.88072504278, 
    1272.68279935669, 
    1262.86251738562, 
    1457.74539290986, 
    1517.71084989314, 
    1728.35885735426, 
    1846.03749934142, 
    1844.66610969961, 
    2159.4268049389, 
    2151.59486453154, 
    2311.2091708874, 
    2441.56767986424, 
    2540.92889054396, 
    2622.28798237923, 
    2701.33265101043, 
    2734.00800824659, 
    2848.60486242213, 
    2912.05264688157, 
    2909.3565168894, 
    2958.22398327703, 
    2922.73579030088, 
    2994.27983055763, 
    3041.84298895705, 
    3045.45367996929, 
    3024.02123351572, 
    2977.17416850313, 
    2875.63941400072, 
    2760.01631381322, 
    2748.70474592129, 
    2661.62403254903, 
    2654.88881668021, 
    2525.295205462, 
    2458.17208878042, 
    2445.35061196372, 
    2456.55232527683, 
    2529.80009173143, 
    2560.32417972254, 
    2694.33413202715, 
    2325.65852594551, 
    2251.01918796174, 
    2106.88810620579, 
    2044.32627043403, 
    1807.15672402228, 
    1576.73053340478, 
    449.057896437575, 
    0, 
    0, 
    0, 
    1143.89708697809, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1023.22406659284, 
    1028.07046624322, 
    858.432058164019, 
    1069.81612445797, 
    1159.10828627412, 
    1481.98055229046, 
    1647.4208814943, 
    1534.10801043554, 
    1798.07827805419, 
    2091.46780137574, 
    2066.60189430994, 
    2170.77277266133, 
    2368.61639021277, 
    2487.16049614065, 
    2493.10870475635, 
    2558.9741485974, 
    2669.18885256918, 
    2717.41825413502, 
    2816.15172327994, 
    2864.10933922811, 
    2813.83580717268, 
    2868.00676993821, 
    3024.25674049923, 
    2877.16429786438, 
    2981.14646377071, 
    3002.46236578491, 
    3027.65716475781, 
    2983.73791272346, 
    2951.29918623495, 
    2903.56137271395, 
    2846.10373104926, 
    2773.44194176221, 
    2668.79210136245, 
    2595.17153502859, 
    2554.92038266444, 
    2452.0963245096, 
    2439.52210758661, 
    2390.92671200997, 
    2480.25951369427, 
    2270.44947082926, 
    2593.12564183396, 
    2484.29355007696, 
    2125.74625293076, 
    2045.98099921541, 
    1900.118571226, 
    1357.28205248142, 
    1027.97071864897, 
    795.46752602101, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1048.14445236103, 
    1146.42211934928, 
    1085.36174487263, 
    1242.62618263092, 
    1346.00374264723, 
    1494.86638579378, 
    1686.7868243678, 
    1843.25368555747, 
    1883.55776665086, 
    2014.99458898156, 
    2076.31280098083, 
    2199.10881326242, 
    2366.25839341113, 
    2447.1236823855, 
    2438.88889674737, 
    2540.85588784398, 
    2645.12654366178, 
    2718.42951326501, 
    2797.51298302309, 
    2843.10584377372, 
    2866.97754763886, 
    3004.86146131239, 
    2887.22732546426, 
    2872.94616678872, 
    2910.22163037332, 
    2955.99707266427, 
    2973.88145882278, 
    2962.6935016814, 
    2936.51658670687, 
    2903.95403774513, 
    2835.61225088129, 
    2766.92410556325, 
    2684.86627654984, 
    2574.12588146134, 
    2536.99155300935, 
    2438.95908758617, 
    2314.81243188305, 
    2216.03624507538, 
    2279.04896540661, 
    2417.58222491708, 
    2274.67708070587, 
    2499.93066435234, 
    2245.9236005366, 
    1921.82698602509, 
    1771.79763879841, 
    1312.75670838663, 
    884.513538089176, 
    630.07914732975, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    960.482809268924, 
    824.718767145798, 
    1078.66930088783, 
    594.375018409947, 
    839.481288223767, 
    1334.06252197331, 
    1412.4707783461, 
    1473.78014044028, 
    1462.11048818373, 
    1545.95237071259, 
    1776.8760268118, 
    1993.53849175443, 
    1976.59805124554, 
    2009.64836108515, 
    2212.26413144658, 
    2357.97378101468, 
    2418.68694274225, 
    2433.59306560811, 
    2522.10617530562, 
    2696.87043523908, 
    2748.05401985648, 
    2821.6295795192, 
    2953.20304589567, 
    2896.69380601961, 
    2859.75285374854, 
    2831.01468086569, 
    2876.12378180113, 
    2917.28119981418, 
    2921.80383421701, 
    2920.57683489112, 
    2911.27184810378, 
    2874.0384647094, 
    2853.34027701088, 
    2799.41323589846, 
    2758.07557007078, 
    2717.29122040693, 
    2676.65178449761, 
    2485.75037031322, 
    2570.2978722836, 
    2390.30346355703, 
    2206.87294147626, 
    2148.9345515403, 
    2160.47027792119, 
    2154.95734317166, 
    2107.15726373147, 
    2246.16371427437, 
    2110.91749435031, 
    1948.1407742292, 
    1626.05329197531, 
    1307.10238961038, 
    573.3402188355, 
    0, 
    0, 
    1199.00615168759, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    919.07793421171, 
    892.324960631045, 
    0, 
    1004.36657910044, 
    838.077694048614, 
    762.285796795296, 
    1164.87034971197, 
    1119.78725919262, 
    1323.63855117028, 
    1641.91015047153, 
    1613.15160501225, 
    1684.55437977202, 
    1862.95324977468, 
    2088.3636470008, 
    2150.70325053416, 
    2114.29910965353, 
    2215.42984982097, 
    2344.18691202434, 
    2364.61856899772, 
    2527.56345332746, 
    2597.33867913488, 
    2682.5608669344, 
    2726.47778735505, 
    2829.67128718485, 
    2827.50561270989, 
    2869.60529253095, 
    2891.35678052611, 
    2885.16610584036, 
    2861.53112699378, 
    2905.145161588, 
    2879.40856566186, 
    2870.96447761723, 
    2845.50695385341, 
    2834.52307818133, 
    2767.56595300677, 
    2763.92304374963, 
    2731.89299001071, 
    2716.33756690141, 
    2703.53092066875, 
    2690.75733388485, 
    2657.25216182512, 
    2487.62309933697, 
    2284.08108601885, 
    2177.11256321605, 
    2059.24054010429, 
    2084.47885033868, 
    2223.06382204398, 
    1975.01887382295, 
    1863.35528412115, 
    2042.49362145299, 
    1836.84692336996, 
    1704.54787616256, 
    1270.88055587705, 
    835.41258449919, 
    1222.35903371197, 
    1440.72812903231, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    498.1099457995, 
    927.81791882338, 
    775.917518537202, 
    840.120187422291, 
    797.060316404972, 
    730.750787504051, 
    917.975335023696, 
    1056.83382000585, 
    1346.7586583238, 
    1373.94225617354, 
    1421.69653628745, 
    1572.84365816086, 
    1707.75305869649, 
    1853.32884326545, 
    1988.607540411, 
    2125.61091906687, 
    2197.25828340569, 
    2209.31128279579, 
    2241.49044108415, 
    2344.56394913092, 
    2463.81830008904, 
    2536.64532513756, 
    2600.25869981975, 
    2691.21392819014, 
    2732.71880364603, 
    2818.29741189643, 
    2818.83101926388, 
    2852.18542368843, 
    2894.97395339196, 
    2892.27505268594, 
    2996.34624437635, 
    2932.23824776554, 
    2884.95319506456, 
    2939.73339309875, 
    2881.71294217081, 
    2927.75130523864, 
    2771.92868700896, 
    2753.07537867922, 
    2677.43613651088, 
    2680.13052983159, 
    2672.49102134569, 
    2696.06063741342, 
    2728.8142524088, 
    2569.55881570843, 
    2396.99984128437, 
    2126.20699092472, 
    2024.08760276637, 
    2038.74637188031, 
    2093.3080075313, 
    1877.58298432554, 
    1920.95238887651, 
    2025.70026737857, 
    1645.75277627852, 
    1818.28055263291, 
    1354.29863537107, 
    1332.60282472167, 
    1663.84708844225, 
    1398.25581649475, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    662.152797667307, 
    840.048587512573, 
    1269.05642106711, 
    872.093470606595, 
    889.097087234037, 
    1231.88562328875, 
    1185.52785160642, 
    1343.87173327895, 
    1483.68725544789, 
    1538.3161078189, 
    1612.05792553987, 
    1806.81167449059, 
    1986.99976832708, 
    2078.7281052802, 
    2233.45133759471, 
    2251.02267652812, 
    2210.11876863801, 
    2263.90703548701, 
    2355.03653294596, 
    2462.92330975131, 
    2545.5159035782, 
    2585.520684178, 
    2661.93784114306, 
    2707.14534943713, 
    2772.80096401747, 
    2833.73151986922, 
    2784.194559859, 
    2768.82346897258, 
    2843.08439094748, 
    2853.41912396534, 
    2806.46353953733, 
    2763.7702973385, 
    2778.59407778709, 
    2787.34555890106, 
    2875.77083051991, 
    2814.4567549669, 
    2687.79921311118, 
    2583.71892099042, 
    2669.73982023091, 
    2626.71887236053, 
    2610.27995680402, 
    2590.33716085167, 
    2662.63729656771, 
    2546.77456600673, 
    2191.53525994501, 
    2015.07027234097, 
    1944.95968641006, 
    1961.84707245294, 
    1906.95987385448, 
    1823.62945168552, 
    1766.78207953795, 
    1357.21085681461, 
    1706.94303687253, 
    1473.34014981246, 
    1374.98469345793, 
    1147.4941578586, 
    1157.42329508638, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    811.341711329656, 
    960.078949389482, 
    788.887327741285, 
    865.674177670456, 
    1078.04887288239, 
    1107.87224004827, 
    1264.38710357394, 
    1376.90490277891, 
    1460.20269877626, 
    1597.38804546017, 
    1639.1244936235, 
    1880.90704318074, 
    2096.21154206596, 
    2215.4691101263, 
    2207.89031829836, 
    2171.09764770011, 
    2188.11159252787, 
    2241.94508527619, 
    2313.59437799983, 
    2412.35032843843, 
    2521.36899579785, 
    2568.36660145256, 
    2631.85652897276, 
    2714.76583058393, 
    2774.5697278596, 
    2797.96786186612, 
    2781.29980330699, 
    2786.67621379463, 
    2837.18049048205, 
    2781.26811291851, 
    2729.2310578574, 
    2763.10595569239, 
    2767.96772562624, 
    2778.62644825491, 
    2806.92451211071, 
    2746.32027238392, 
    2621.10304063611, 
    2566.29293252912, 
    2535.28280784861, 
    2607.27143770612, 
    2527.4877069102, 
    2480.95759649024, 
    2514.79816997184, 
    2445.84574128953, 
    2207.12858811114, 
    1992.79354621248, 
    1896.58045398186, 
    1908.99898239662, 
    1748.31241812206, 
    1920.17161462801, 
    1670.15764715738, 
    1626.34306856918, 
    1691.67611803836, 
    1098.63741155899, 
    827.84326837381, 
    789.246383328462, 
    964.553290037875, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    1011.23560833829, 
    1053.51467246011, 
    849.980323179244, 
    851.986281398676, 
    936.278712141493, 
    1158.84339050702, 
    1201.26927576888, 
    1294.14088774858, 
    1441.35201531952, 
    1605.02950305208, 
    1632.38653892047, 
    1900.82925905572, 
    2120.02044941242, 
    2140.82210488796, 
    2003.23597927256, 
    2029.90930705656, 
    2145.97784326414, 
    2260.46962604304, 
    2322.11623106821, 
    2375.38531278005, 
    2488.51199324252, 
    2547.65447652582, 
    2592.47128137274, 
    2604.57862750184, 
    2711.99951029191, 
    2767.42137352793, 
    2795.34790374321, 
    2737.04939536208, 
    2741.47783871447, 
    2717.62978040104, 
    2684.99542473884, 
    2726.10021739774, 
    2723.80552882712, 
    2658.15882510747, 
    2605.49601111018, 
    2547.29852537951, 
    2575.41226642714, 
    2564.58252438774, 
    2517.41906319918, 
    2578.47352370503, 
    2449.76587695291, 
    2379.20574079118, 
    2354.70904643882, 
    2345.86998046125, 
    2233.44662606884, 
    2093.41724425281, 
    1900.84003285931, 
    1925.0748435489, 
    1873.77840744428, 
    2039.64468801157, 
    2004.91219058222, 
    1786.26308920577, 
    1350.31278820692, 
    1003.61689311722, 
    795.222096101771, 
    757.391477234823, 
    988.696342767115, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    223.781026122609, 
    471.835215462414, 
    667.362675750979, 
    616.416974442618, 
    838.019606433519, 
    940.233916107683, 
    1059.38304734698, 
    1235.18890440776, 
    1260.25002213328, 
    1438.66835294796, 
    1539.62493691843, 
    1635.65956894162, 
    1901.50076285264, 
    1993.03675602844, 
    1821.0200774261, 
    1913.50757572026, 
    2068.48035139895, 
    2142.26570929789, 
    2226.73618411146, 
    2272.58477204943, 
    2366.84788561199, 
    2501.09971996401, 
    2504.67765347737, 
    2544.44127953989, 
    2563.49161066965, 
    2625.45971269977, 
    2703.15319361072, 
    2808.29527671875, 
    2726.83509861083, 
    2725.77803132008, 
    2715.54384129582, 
    2688.84436484561, 
    2723.26780957174, 
    2715.83049625054, 
    2612.71642765592, 
    2679.85217154967, 
    2630.65929595966, 
    2621.86927651957, 
    2558.91788286748, 
    2490.70237379423, 
    2420.38053191544, 
    2357.89678723107, 
    2292.21308040672, 
    2282.30352138107, 
    2297.35042295652, 
    2188.89435547139, 
    2212.07405270254, 
    1873.58067317311, 
    1763.17624912184, 
    1737.10965346444, 
    1877.01560683459, 
    2037.36660268074, 
    2002.36089556024, 
    1520.56654386129, 
    770.512013559677, 
    972.629452917414, 
    731.074721387138, 
    170.665849463938, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    783.298286077705, 
    734.775851623196, 
    1414.7179092718, 
    1296.37800375321, 
    1396.376048336, 
    1492.6074695572, 
    1656.9662708266, 
    1883.84154977545, 
    1787.59991326103, 
    1733.98025995536, 
    1885.87780814727, 
    2014.11723345116, 
    2102.036036793, 
    2196.29069474978, 
    2272.86854542233, 
    2326.94361656102, 
    2418.59257087225, 
    2432.76600582868, 
    2473.46851411382, 
    2511.99044582416, 
    2579.51851881891, 
    2604.2883915771, 
    2655.67903755951, 
    2664.82592307674, 
    2721.77828311319, 
    2721.70161522425, 
    2676.06084981524, 
    2701.73527935093, 
    2722.63547026402, 
    2565.60209880457, 
    2569.44378749146, 
    2543.05164612605, 
    2548.25183363521, 
    2437.94378647697, 
    2391.64514867424, 
    2350.66780992792, 
    2303.85093529254, 
    2278.98268799178, 
    2268.49618353863, 
    2275.35869074778, 
    2111.85778931155, 
    1954.50099148355, 
    1992.74982127288, 
    1826.52082981262, 
    1807.45037123165, 
    1941.70325203798, 
    2073.73931917488, 
    2069.41165583263, 
    1655.58259035695, 
    1022.56321971504, 
    1153.89802118759, 
    1021.43213908258, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1031.65018623117, 
    1384.82772100866, 
    1218.42886884058, 
    1283.35460061752, 
    1431.92912853956, 
    1566.99665187902, 
    1683.77722397336, 
    1652.23739044544, 
    1761.01017756568, 
    2007.65290059248, 
    2049.92839554524, 
    2042.5556045387, 
    2133.08505618563, 
    2230.41434160296, 
    2331.72521141869, 
    2324.84208188489, 
    2385.57266758091, 
    2483.4671223021, 
    2485.61091661573, 
    2534.45557589996, 
    2524.25739084788, 
    2511.68606847295, 
    2578.86640075547, 
    2681.4829705531, 
    2699.89403293438, 
    2647.33141621615, 
    2671.63641630283, 
    2645.21414193042, 
    2574.11465398235, 
    2547.92913426725, 
    2501.71643293117, 
    2512.33843705306, 
    2419.73621066947, 
    2370.64813628373, 
    2351.65414533204, 
    2304.1202934805, 
    2255.36900918779, 
    2209.32546339301, 
    2109.68811751072, 
    1934.12318723305, 
    1973.53218507677, 
    1936.91264329023, 
    1785.53186181735, 
    1779.81333904695, 
    1594.08290657658, 
    1951.67807788466, 
    2048.21765294452, 
    1705.36495179627, 
    807.893889942032, 
    755.573958661416, 
    1134.34880674418, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    656.379692004648, 
    900.481277762625, 
    851.801287595232, 
    1073.46505440119, 
    1203.29760154092, 
    1345.97082870116, 
    1365.47899460939, 
    1424.61428901853, 
    1515.29490207206, 
    1580.37751128538, 
    1721.63341030731, 
    1919.72387080464, 
    1907.81666838407, 
    1968.10730925134, 
    2087.74761820109, 
    2148.30602528012, 
    2232.07995014398, 
    2264.87846705772, 
    2359.84467112148, 
    2506.8289339751, 
    2480.50433588607, 
    2497.70992399396, 
    2461.68772676835, 
    2488.72592359834, 
    2523.80209327368, 
    2630.90654465522, 
    2638.71516557238, 
    2637.92098709148, 
    2622.53735185866, 
    2600.78196918484, 
    2572.79945394804, 
    2539.11548173781, 
    2572.93603895274, 
    2539.10774994575, 
    2408.100496263, 
    2365.31187443165, 
    2368.99060610861, 
    2297.77900122195, 
    2217.14192364782, 
    2157.67058566652, 
    1999.64301475306, 
    1896.66942075434, 
    1891.94305253428, 
    1884.81220810037, 
    1758.58874499482, 
    1833.06105164243, 
    1807.94511095742, 
    2011.43678433413, 
    2069.79970796433, 
    1706.02439791699, 
    1024.98451741513, 
    743.280046099653, 
    750.80421908493, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    795.925864718975, 
    643.099088259866, 
    919.48541972384, 
    1024.39812559998, 
    1180.2801919529, 
    1212.4007733735, 
    1271.82088087861, 
    1343.19667537998, 
    1396.25905024119, 
    1491.26910771014, 
    1644.46643674319, 
    1800.88739618778, 
    1815.17628293971, 
    1904.24240089446, 
    2064.80241712352, 
    2115.44843582758, 
    2127.14345558638, 
    2276.73102732051, 
    2388.53738866801, 
    2383.42619003635, 
    2426.63047276119, 
    2414.50387239872, 
    2413.08593912344, 
    2435.82024348265, 
    2464.48120532147, 
    2574.78181030699, 
    2535.30206411195, 
    2552.60439771631, 
    2547.55360950638, 
    2548.73946052931, 
    2513.73271194526, 
    2506.65409030136, 
    2418.27610864217, 
    2452.19803868251, 
    2407.44438778353, 
    2375.45894970108, 
    2312.57645865077, 
    2251.41486041008, 
    2168.05540596459, 
    2012.55147757653, 
    1921.08216119123, 
    1851.98862928521, 
    1860.40125862273, 
    1841.92727118192, 
    1806.97528455347, 
    1788.47248288766, 
    1884.20264359516, 
    1887.28697191938, 
    1936.58038535303, 
    1819.91662798049, 
    1488.06424392484, 
    1348.59979488066, 
    1072.75875079461, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    813.284107287358, 
    759.46610706028, 
    927.897916349777, 
    1020.8503363388, 
    1028.17596588818, 
    1111.3312533981, 
    1205.53910902048, 
    1165.58957761291, 
    1244.44727977178, 
    1349.71973339045, 
    1447.3086669056, 
    1591.21584526624, 
    1731.85195036404, 
    1832.11541505061, 
    1854.23425464497, 
    1932.44854014731, 
    2077.49030892287, 
    2070.70577002865, 
    2179.90849969922, 
    2235.33983469609, 
    2306.31134492534, 
    2331.89875847642, 
    2310.94543181837, 
    2294.37854937529, 
    2451.16732499805, 
    2430.02807734446, 
    2439.74103599027, 
    2448.53001021774, 
    2437.50727038209, 
    2495.34677666049, 
    2525.12349182594, 
    2495.02252454181, 
    2496.55231557723, 
    2428.72639711729, 
    2404.51421042335, 
    2368.01062612215, 
    2372.37099270417, 
    2256.31460665896, 
    2210.4418496899, 
    2159.79745799241, 
    1995.64796649074, 
    1883.14394118453, 
    1827.35998348247, 
    1827.66264687381, 
    1748.63265336495, 
    1682.6256221483, 
    1794.14689916417, 
    1901.90843628551, 
    1803.04723554234, 
    1814.08379053388, 
    1721.22014997943, 
    1700.08109124393, 
    1666.74794655743, 
    1559.25086844357, 
    1040.7855418629, 
    101.642078103247, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    736.695486954855, 
    887.007338573262, 
    942.990916512837, 
    877.906482366629, 
    889.530596701368, 
    951.969724621112, 
    962.474558111996, 
    1076.42740060409, 
    1053.23891337996, 
    1140.99981319223, 
    1287.7600617861, 
    1397.27172132101, 
    1521.26066927106, 
    1669.24358481948, 
    1758.5916974566, 
    1773.30572341929, 
    1902.96468562737, 
    1972.9481859751, 
    2016.39340506957, 
    2062.48061111947, 
    2140.1932340076, 
    2199.88385665783, 
    2207.42661023957, 
    2234.09692089187, 
    2181.06219832937, 
    2516.73923627286, 
    2323.86691731978, 
    2298.49739299744, 
    2312.06234309858, 
    2311.64045703575, 
    2307.73996846131, 
    2409.73703887806, 
    2472.22511372819, 
    2459.87623895451, 
    2368.86786508147, 
    2317.7635365702, 
    2351.49703364568, 
    2279.50372173745, 
    2252.38091354117, 
    2172.66692254124, 
    2096.14307857633, 
    1991.40688211688, 
    1855.0593683105, 
    1789.43131040621, 
    1758.15700325325, 
    1731.73076009394, 
    1755.24158164107, 
    1775.84192921446, 
    1785.05666911498, 
    1669.97515287504, 
    1609.34160743064, 
    1650.40423756612, 
    1571.44729108299, 
    1015.70855298054, 
    563.231741625589, 
    869.921334330832, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    867.740232559925, 
    682.063689926776, 
    679.809120971515, 
    737.793317807865, 
    668.159458177931, 
    0, 
    689.280152169446, 
    974.249955143302, 
    898.499168587703, 
    928.122975190973, 
    1068.12667962498, 
    1190.01416840563, 
    1329.38712507131, 
    1460.78067813321, 
    1594.02484936203, 
    1664.81621907929, 
    1803.91506565592, 
    1838.19649085969, 
    1909.0126067735, 
    1942.05125145653, 
    1992.18205511138, 
    2038.29555831788, 
    2104.70882369636, 
    2124.19803304195, 
    2120.77479374581, 
    2099.12376200139, 
    2463.68126483905, 
    2111.25103078079, 
    2231.33185823434, 
    2269.81401303126, 
    2223.38395470542, 
    2203.90328531221, 
    2316.21984938176, 
    2414.08842000847, 
    2387.71207328327, 
    2312.7739358739, 
    2218.0794029261, 
    2204.0904299797, 
    2192.38151859469, 
    2135.49552597536, 
    2059.05757803275, 
    1986.46206649726, 
    1910.02600755009, 
    1787.86433121661, 
    1679.94667500241, 
    1605.23830323098, 
    1559.5395341819, 
    1589.89478208244, 
    1617.35453557168, 
    1638.30458480916, 
    1468.27743867978, 
    1344.65189741454, 
    1472.3765724008, 
    1755.69193155439, 
    328.604994633085, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    695.654112776919, 
    402.258887223841, 
    652.852166712489, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1046.7501589799, 
    816.206050274473, 
    1068.3937129759, 
    1156.90215849313, 
    1297.33599341501, 
    1438.80735039763, 
    1540.98957808229, 
    1637.07385321361, 
    1698.6773062008, 
    1758.21820005247, 
    1812.66319961529, 
    1894.00496720145, 
    1951.38049761256, 
    1945.39155130003, 
    2006.65426771846, 
    2025.06961837396, 
    1999.8243816096, 
    1939.36073151536, 
    2309.0385652095, 
    2156.1042362757, 
    2203.85003691239, 
    2242.4442707392, 
    2155.54393737349, 
    2239.71100766276, 
    2260.81814306991, 
    2332.98048311914, 
    2370.58963652205, 
    2265.59411736655, 
    2060.67636451273, 
    2016.09253472054, 
    2114.9078648471, 
    2040.21148772893, 
    2018.33825268525, 
    1949.67597468841, 
    1817.20032788949, 
    1701.83389899775, 
    1595.76516336986, 
    1473.20029571043, 
    1355.64397060001, 
    1346.8146988798, 
    1292.54720287474, 
    1476.6618597255, 
    1383.88677666714, 
    1193.41894558605, 
    1166.20877890383, 
    1259.9625440217, 
    1299.81389508319, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    768.330592171638, 
    1055.69682430308, 
    1177.23464705179, 
    1274.88198824948, 
    1447.08012666015, 
    1521.31661631907, 
    1557.1360857014, 
    1618.11870945145, 
    1555.7900358979, 
    1757.1949891895, 
    1857.1272864178, 
    1964.41921048815, 
    1961.56188698752, 
    1917.79623568595, 
    1925.64063356081, 
    1915.61947108333, 
    1937.48544542606, 
    2268.64356902712, 
    2073.2637081319, 
    2137.35058405793, 
    2215.21629134044, 
    2191.51434328129, 
    2191.60363519464, 
    2124.49430610581, 
    2246.21797859668, 
    2253.29620974711, 
    2272.86623139094, 
    2090.20604217965, 
    1944.27401346881, 
    2041.245523587, 
    2104.74440601348, 
    2009.391385099, 
    1875.24658628465, 
    1755.24898453194, 
    1633.57025841454, 
    1517.10114262154, 
    1385.46232955659, 
    1250.00839323954, 
    1163.57627070883, 
    1098.40395284601, 
    1454.4061509468, 
    1201.70595812631, 
    859.808051735083, 
    737.536573564025, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    840.171609686753, 
    1125.02403064185, 
    1100.7554190044, 
    1176.57074889457, 
    1347.45662912852, 
    1424.69844431936, 
    1498.75848529854, 
    1506.95324821699, 
    1324.29301771533, 
    1407.65197995495, 
    1710.04056720828, 
    1849.83622745897, 
    1966.06911245152, 
    2085.99625448698, 
    2012.47058933823, 
    1942.44842612542, 
    1945.15996097574, 
    2168.39506097609, 
    1962.89515214844, 
    1958.96477094651, 
    2048.73068532145, 
    2005.1086867454, 
    1977.2865162881, 
    2093.61533380711, 
    2086.31745434806, 
    2053.92664564909, 
    1984.5774835388, 
    2159.34746295263, 
    2114.12121280702, 
    1815.17818473886, 
    1985.83603483512, 
    1997.11826855323, 
    1958.60687905462, 
    1814.71650100856, 
    1672.00518224402, 
    1542.84651195648, 
    1434.97078809293, 
    1197.99903090775, 
    1193.65640381984, 
    1076.90509341726, 
    1098.14045666416, 
    1126.08440058995, 
    828.355785621388, 
    872.436734778291, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1108.77164591924, 
    1321.87671223413, 
    1452.30642294477, 
    1461.63730692852, 
    1092.19279310866, 
    947.900085304985, 
    1291.38487602415, 
    1534.22245987956, 
    1844.81890018964, 
    2018.28338260949, 
    2033.36492443385, 
    1888.31537650252, 
    1701.92790688495, 
    1963.66009262491, 
    1784.97600621501, 
    1744.6313161633, 
    1952.59910675545, 
    1942.30908237073, 
    1700.08167466184, 
    1769.9453850284, 
    1947.60305751998, 
    1903.189889761, 
    1920.0982475706, 
    1896.34955496475, 
    2040.56649119293, 
    1984.95736154053, 
    1920.46735476067, 
    2028.92250590045, 
    2025.09779679143, 
    1919.54124522959, 
    1759.90388622121, 
    1554.06767328467, 
    1404.96612392705, 
    1352.50989726964, 
    1139.65252221837, 
    880.013639141899, 
    1083.65546506142, 
    900.576990513901, 
    1107.8969923275, 
    845.2606887542, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1171.20899442683, 
    1203.12171867719, 
    1174.94968664839, 
    722.725131184243, 
    839.769374600437, 
    899.177670458785, 
    1022.63344620995, 
    1695.12434136002, 
    1897.98928753515, 
    1791.00304368405, 
    1710.98450462882, 
    1720.55388902982, 
    1713.09877812453, 
    1766.89529132947, 
    1637.43038568638, 
    1542.91112329001, 
    1583.19570515741, 
    1734.06245984595, 
    1670.98066912761, 
    1773.74920233509, 
    1702.85864398471, 
    1730.22502266448, 
    1699.74017809079, 
    1797.40245638125, 
    1930.16925506078, 
    1761.18513429965, 
    1832.21934096391, 
    1868.0168808876, 
    1902.68187074951, 
    1870.85016606676, 
    1643.6236150195, 
    1439.4589088969, 
    1263.99587891753, 
    1090.54795852381, 
    902.014386691376, 
    789.575042691679, 
    838.615748698646, 
    43.3933025530239, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    822.205957761807, 
    1230.07024100286, 
    1938.53456627146, 
    1880.55103179938, 
    1455.07564550387, 
    1342.20016237123, 
    1449.78519853645, 
    1627.83939136447, 
    1724.73207089323, 
    1453.16856025111, 
    1435.24399262452, 
    1663.13300092243, 
    1551.79621911613, 
    1622.67286580426, 
    1504.73694398318, 
    1573.56695727707, 
    1660.1897069044, 
    1531.40912763024, 
    1615.09339068712, 
    1679.16494193395, 
    1581.25105530098, 
    1637.37700414338, 
    1503.21090656994, 
    1497.43138470633, 
    1653.12531102964, 
    1754.81810867173, 
    1501.582948592, 
    1215.21620821175, 
    1041.95571999276, 
    808.748032788677, 
    618.964278506231, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    909.455874871708, 
    1503.7903722337, 
    1665.59424751957, 
    1245.36657857209, 
    1232.57954912647, 
    1353.11436433668, 
    1424.47652659997, 
    1382.00540442789, 
    1613.31567090478, 
    1260.61442955182, 
    1385.86870177165, 
    1629.41533983879, 
    1752.23195092564, 
    1363.04110533616, 
    1315.33468045601, 
    1513.60439574335, 
    1583.08788836968, 
    1492.93651120653, 
    1469.42713487761, 
    1500.47653653459, 
    1475.79708573943, 
    1362.80767442505, 
    1409.90751409869, 
    1355.04513840894, 
    1372.31994497558, 
    1632.73146764407, 
    1580.41884239273, 
    1319.66303528665, 
    972.364941408943, 
    780.991248877619, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    741.451375949156, 
    1374.72472608478, 
    964.889104021041, 
    1227.92219993612, 
    1210.65978957111, 
    1152.88734282373, 
    1099.01811787837, 
    1169.58882727002, 
    1375.44495713084, 
    1156.13649549529, 
    1241.24612065519, 
    2001.00816759498, 
    1417.28097355999, 
    1293.96497799644, 
    1121.25030572989, 
    1317.06974833328, 
    1357.21784266745, 
    1210.71332427556, 
    1360.35897832401, 
    1442.74324959804, 
    1328.58495034445, 
    1234.67273814119, 
    1359.22387105718, 
    1142.9787830832, 
    1043.74750630126, 
    1458.88092475789, 
    1645.36955928121, 
    960.448118514539, 
    1276.56655537612, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    529.585423514496, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1174.30608227374, 
    760.11972141423, 
    818.679343580324, 
    1047.81895005274, 
    803.398676595915, 
    727.849023224591, 
    942.435989465244, 
    916.632130160548, 
    937.203173225275, 
    920.079268155583, 
    1652.08982560871, 
    1055.42868426198, 
    1050.12964629921, 
    1034.52452792101, 
    1322.71826600555, 
    1165.6706267914, 
    868.859422289162, 
    1021.88021429658, 
    1219.34178215208, 
    1171.22675984497, 
    1139.63308708865, 
    1158.85575614324, 
    923.256625927131, 
    1076.27350464859, 
    1215.93435924992, 
    908.904313195504, 
    0, 
    869.801224874338, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    573.713421166239, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1012.15339859553, 
    834.761038951223, 
    781.22917100357, 
    0, 
    0, 
    934.177099524366, 
    0, 
    1046.44942598694, 
    1611.51987857977, 
    786.123843959548, 
    800.273351827993, 
    1054.04092233291, 
    1557.85101334603, 
    1005.11942528085, 
    781.543803048291, 
    851.939243532074, 
    1020.03984736201, 
    1049.43512193782, 
    998.740183895374, 
    661.068376047252, 
    770.645615196513, 
    0, 
    1098.45003070636, 
    0, 
    0, 
    0, 
    32.3741719330262, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    611.102052959641, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1149.7709516235, 
    0, 
    0, 
    899.345270510427, 
    1118.97260456218, 
    679.594972934562, 
    1058.99306418638, 
    734.077593447327, 
    699.732642440551, 
    782.015681196706, 
    594.730213526081, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    836.536915679264, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    930.577676060031, 
    0, 
    0, 
    0, 
    0, 
    0, 
    733.582189673009, 
    0, 
    0, 
    633.41550416689, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    792.340430466792, 
    629.787205834943, 
    652.420853123232, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    709.311850782452, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    364.860236785387, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0 ;

 topg =
  
    -3407.00706531486, 
    -3447.89348203311, 
    -3469.7266554197, 
    -3473.83785846706, 
    -3441.45892785084, 
    -3455.66498616081, 
    -3427.45636919284, 
    -3419.87941848738, 
    -3395.47319972261, 
    -3326.86166316905, 
    -3313.43655655232, 
    -3260.88644908123, 
    -3194.15038720758, 
    -3100.50494213895, 
    -3023.62121482926, 
    -2848.92162949241, 
    -2784.27391706682, 
    -2405.14896549169, 
    -2292.20102496003, 
    -2195.07834583381, 
    -2045.31040587217, 
    -1951.86944313519, 
    -1639.0241496053, 
    -1485.42673783767, 
    -943.229973471577, 
    -602.13016587756, 
    -518.75648005572, 
    -930.576852633999, 
    -1230.59214360663, 
    -1480.72905186977, 
    -1849.15177015281, 
    -1961.45523035406, 
    -2138.6434976849, 
    -2261.04156979415, 
    -2461.40437930322, 
    -2575.33448386539, 
    -2636.2243837568, 
    -2805.14913947265, 
    -2895.99494153201, 
    -2859.39492780764, 
    -2919.3359911877, 
    -2931.70152810707, 
    -2960.03166456746, 
    -3039.15411793879, 
    -3030.66700390926, 
    -3068.24406250273, 
    -3029.73705408795, 
    -2978.58828605489, 
    -2861.42159111476, 
    -2974.57541272889, 
    -2947.30233716805, 
    -2946.35860426882, 
    -3013.72315908947, 
    -2804.42944841716, 
    -2682.07476878407, 
    -2728.38689457636, 
    -2609.24997095191, 
    -2436.61347447104, 
    -2341.95395037575, 
    -2351.87962818039, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3420.50206774533, 
    -3438.21536196787, 
    -3417.37483500687, 
    -3418.59141774621, 
    -3425.06951378014, 
    -3414.68342557867, 
    -3409.49723052124, 
    -3393.88246966423, 
    -3364.6341143669, 
    -3330.18171854222, 
    -3274.02916694462, 
    -3245.50968873301, 
    -3164.55481507236, 
    -3085.80320184415, 
    -2993.85755689734, 
    -2920.97674440937, 
    -2653.26889342236, 
    -2152.55345237535, 
    -2015.20702766171, 
    -1829.16528532192, 
    -1171.5143949844, 
    -564.201956139163, 
    -285.316292586544, 
    -208.853331457994, 
    -387.57825417855, 
    -182.785081763017, 
    -183.143711871823, 
    -199.427389080821, 
    -316.263631293113, 
    -781.752310074725, 
    -1351.1722069342, 
    -1802.28694123784, 
    -1958.56777755891, 
    -2114.2177778118, 
    -2298.64551358794, 
    -2416.41396954612, 
    -2676.59635810809, 
    -2694.35453863026, 
    -2804.91421505372, 
    -2866.0365347355, 
    -2868.92884660915, 
    -2885.12726581911, 
    -2948.45942788802, 
    -3016.99574701837, 
    -3042.97362956595, 
    -3035.03746386418, 
    -3021.79662228165, 
    -2914.37875366211, 
    -2870.30030205909, 
    -2843.95451373776, 
    -2737.2669487384, 
    -2882.44931009769, 
    -2931.56529131608, 
    -2638.22948497674, 
    -2558.22940596594, 
    -2735.90699745853, 
    -2612.26775880409, 
    -2274.69938821996, 
    -2276.2431791675, 
    -2249.40315839505, 
    -2099.14159062675, 
    -2294.83908562911, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3450.27360912293, 
    -3429.24417445748, 
    -3405.99251912663, 
    -3408.67583404917, 
    -3409.7092361023, 
    -3405.05653663285, 
    -3392.20106719937, 
    -3390.60958383866, 
    -3351.71848668764, 
    -3328.10484995741, 
    -3274.8883062792, 
    -3228.1872942712, 
    -3151.81661734416, 
    -3100.31450206248, 
    -3033.93864473383, 
    -2835.11485534873, 
    -2521.55004482974, 
    -2382.39628250788, 
    -1578.92784484316, 
    -695.369056488069, 
    -200.018697275159, 
    -154.728684511857, 
    -140.821784889845, 
    -149.398396386278, 
    -145.425219865822, 
    -119.808299962777, 
    -116.09636588166, 
    -150.116817106992, 
    -182.032381707049, 
    -195.495610122852, 
    -491.181472146101, 
    -1655.60899775079, 
    -1847.40051609565, 
    -1965.51343145936, 
    -2161.12682500585, 
    -2440.0095686448, 
    -2570.44053238103, 
    -2587.7943339759, 
    -2670.39787574418, 
    -2706.14063135641, 
    -2789.41687807978, 
    -2922.82205251457, 
    -2946.46880809617, 
    -3006.09799290024, 
    -3019.73474876344, 
    -3035.4927097846, 
    -3014.19561859848, 
    -3016.24762871925, 
    -2984.9835803127, 
    -2970.0424804004, 
    -2800.53151184287, 
    -2951.54179155066, 
    -3163.16195603528, 
    -2995.14105826076, 
    -2659.36606668812, 
    -2597.08217341475, 
    -2896.08956300878, 
    -2396.16043675199, 
    -2336.73470532801, 
    -2251.76287072877, 
    -2108.72441637609, 
    -1873.52237107639, 
    -2265.30835972494, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3396.35830425335, 
    -3384.24891534444, 
    -3392.64375296632, 
    -3396.06761909305, 
    -3400.19957645156, 
    -3392.28707858403, 
    -3399.21385638845, 
    -3368.26409020162, 
    -3341.15864363069, 
    -3313.86415197494, 
    -3261.41380509978, 
    -3239.7791971888, 
    -3166.14617947261, 
    -2945.61982417774, 
    -2947.67357175, 
    -2858.53042992125, 
    -2629.21541821863, 
    -2026.70710371643, 
    -1428.25212326135, 
    -247.252603253216, 
    -137.076724587469, 
    -125.510156816224, 
    -113.559198631551, 
    -94.0510473165904, 
    -15.0301875435349, 
    339.807780096009, 
    155.636467769192, 
    7.99177745208328, 
    -116.902752287844, 
    -180.70750452236, 
    -204.398211450353, 
    -1069.45233583183, 
    -1775.80802099008, 
    -1916.40294120079, 
    -2180.90729467172, 
    -2354.18872022469, 
    -2577.9647046951, 
    -2479.45160400801, 
    -2566.02937636423, 
    -2677.89155214658, 
    -2760.07483747425, 
    -2864.59397507141, 
    -2948.54923244019, 
    -2992.09819384465, 
    -2992.36726210232, 
    -3018.77708853693, 
    -2860.23613422048, 
    -2987.06264544548, 
    -2975.22980190845, 
    -2950.35464156301, 
    -2982.92332272247, 
    -3029.10041356274, 
    -3064.43521562429, 
    -2983.1411032682, 
    -2619.29385099165, 
    -2639.77397352264, 
    -2742.07141499449, 
    -2440.06472152932, 
    -2275.14254412165, 
    -2271.83283530104, 
    -2175.77363909372, 
    -1873.30621129428, 
    -1807.41446158654, 
    -2219.41365722793, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3368.74221747079, 
    -3367.14321041641, 
    -3395.48095327209, 
    -3366.76524542694, 
    -3366.99670023988, 
    -3376.70864977522, 
    -3375.39937582155, 
    -3338.43490433132, 
    -3296.79702300854, 
    -3253.38361115151, 
    -3180.61310422754, 
    -3121.42367953549, 
    -3082.00813671082, 
    -2998.25563485038, 
    -2879.07586546895, 
    -2799.32244394608, 
    -2617.93015958267, 
    -1824.9204186998, 
    -750.037060638281, 
    -124.50756300043, 
    -119.392913904863, 
    -88.1948156805342, 
    -1.51972247988865, 
    196.623743941515, 
    272.132601687785, 
    282.413272879026, 
    635.17194914097, 
    489.102854007836, 
    53.0620013475422, 
    -166.575533684264, 
    -195.904899868426, 
    -526.027195532138, 
    -1708.34947245599, 
    -1955.19091195409, 
    -2049.94794434209, 
    -2250.17351618272, 
    -2478.83154590773, 
    -2421.43085916312, 
    -2479.58563543407, 
    -2656.26737865008, 
    -2749.76385405777, 
    -2834.41368210676, 
    -2940.6160797085, 
    -2984.71852373249, 
    -2983.19282239549, 
    -2981.02296907397, 
    -2944.51716133622, 
    -2963.99190115421, 
    -2980.01606335271, 
    -2987.13720836404, 
    -2897.60176300014, 
    -2981.49406417727, 
    -2901.32579479666, 
    -2916.04085972221, 
    -2873.53279645179, 
    -2645.56364709186, 
    -2621.50520972308, 
    -2387.87481832985, 
    -2411.94058138686, 
    -2290.62319983881, 
    -2248.29443574673, 
    -2010.75247371797, 
    -1871.26153617423, 
    -1731.21898265809, 
    -2008.28201830481, 
    -2299.33070211208, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3384.05609568289, 
    -3380.45029332416, 
    -3357.50817782241, 
    -3348.08436032559, 
    -3349.1613362858, 
    -3366.70343817255, 
    -3337.60193838224, 
    -3277.45276917802, 
    -3213.19549270066, 
    -3149.30715487866, 
    -3076.34647867474, 
    -2990.68892000717, 
    -2926.19003617136, 
    -2987.3838351977, 
    -2833.83906163881, 
    -2550.95893502742, 
    -1336.65818776368, 
    -1392.32679259843, 
    -540.051676836687, 
    -105.97666677302, 
    -89.6844285685163, 
    -61.8723504343063, 
    99.5245890110104, 
    192.503628153017, 
    934.015541845575, 
    584.424185407928, 
    1012.99867482628, 
    910.089751744454, 
    211.555196696141, 
    -205.430450665858, 
    -335.067964850726, 
    -386.578121753448, 
    -1355.17543265588, 
    -1772.61272176676, 
    -1848.15708350921, 
    -1984.71444584248, 
    -2279.85476294985, 
    -2446.83330287271, 
    -2548.06478294039, 
    -2703.05824438695, 
    -2775.68375775208, 
    -2865.86096656176, 
    -2920.64990258297, 
    -2922.84952786949, 
    -2961.21259430034, 
    -2996.09944660319, 
    -2985.37247189375, 
    -2979.52636394095, 
    -2975.63386841504, 
    -2979.04931910601, 
    -2878.52714591544, 
    -2973.03388250849, 
    -2978.60379957859, 
    -2948.05959980485, 
    -2843.39099206529, 
    -2808.31029313142, 
    -2733.36756331389, 
    -2474.76471104467, 
    -2391.93215344334, 
    -2320.44541772242, 
    -2282.12575894107, 
    -2133.69590535436, 
    -1833.5357440124, 
    -1736.22882074952, 
    -1632.28885343921, 
    -1684.18650026738, 
    -2299.04662047041, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3328.40387612201, 
    -3327.12849742381, 
    -3317.23964346857, 
    -3322.22589176259, 
    -3315.53086694117, 
    -3277.62891742497, 
    -3225.22985378492, 
    -3167.053489967, 
    -3119.56413937149, 
    -3052.29409595246, 
    -3026.62398875067, 
    -2897.47155806145, 
    -2824.84613549723, 
    -2733.14854873708, 
    -2455.33256693088, 
    -728.712438547052, 
    -212.932035555095, 
    -413.169254785691, 
    -199.909659677233, 
    -117.439683991077, 
    -93.3678447012138, 
    -27.4592920720635, 
    300.023374512634, 
    414.229781916534, 
    584.98605373165, 
    1057.4383658722, 
    810.874473956234, 
    750.155046050783, 
    -13.4711116526978, 
    -106.033484844451, 
    -215.001901009315, 
    -185.749713923336, 
    -1201.93068226028, 
    -1741.7331759975, 
    -1953.36770394081, 
    -2076.77646229436, 
    -2431.1778196055, 
    -2478.96767012883, 
    -2563.41074124429, 
    -2662.98959207054, 
    -2799.39766167687, 
    -2856.00619028397, 
    -2894.87457138694, 
    -2890.1286699011, 
    -2917.21705434357, 
    -2918.83684755947, 
    -2924.18739200947, 
    -2933.31538813165, 
    -2924.77173330002, 
    -2975.03370637456, 
    -2898.23082508459, 
    -2931.60569450489, 
    -2801.61335287916, 
    -2718.84114640291, 
    -2733.5071512972, 
    -2817.71604001855, 
    -2743.02475344667, 
    -2498.77434814043, 
    -2433.62215858451, 
    -2379.12066667478, 
    -2251.71766243964, 
    -2216.02808416864, 
    -2027.30420258491, 
    -1871.85404494949, 
    -1684.28263198835, 
    -1591.85788789174, 
    -1539.66819698252, 
    -2280.11536878221, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3304.7544264158, 
    -3300.91566397228, 
    -3296.5194796811, 
    -3295.79424392683, 
    -3280.74079479803, 
    -3223.34510473441, 
    -3156.01874264571, 
    -3093.9072395487, 
    -3015.50315643345, 
    -2955.76309528757, 
    -2892.12110810317, 
    -2855.51751606462, 
    -2721.47134648886, 
    -1675.8861949959, 
    -187.647010053523, 
    -120.558232546654, 
    -108.483513871606, 
    -458.891541082676, 
    -352.123665936714, 
    -156.634210556648, 
    -12.1294357801998, 
    107.572358445387, 
    167.869721230577, 
    642.443841248589, 
    713.728226536732, 
    1019.20060025991, 
    725.983245460898, 
    541.734606632869, 
    471.228603038381, 
    137.96989430479, 
    -219.161078202099, 
    -404.628322878988, 
    -724.588015950411, 
    -1762.21096080682, 
    -1990.26432897689, 
    -2032.40006815706, 
    -2333.24502020106, 
    -2347.76035837684, 
    -2484.83660434155, 
    -2617.34899909179, 
    -2702.01713413354, 
    -2815.58772446994, 
    -2874.97413346482, 
    -2888.10212377738, 
    -2882.01794474603, 
    -2899.29459749331, 
    -2895.14268160454, 
    -2910.9260111058, 
    -2913.98100255131, 
    -2918.73263802694, 
    -2933.23830267724, 
    -2932.70589868219, 
    -2880.6459689936, 
    -2834.11864209149, 
    -2840.37040664314, 
    -2664.67759501253, 
    -2758.81862589974, 
    -2561.8618241638, 
    -2499.01925583996, 
    -2417.79919806093, 
    -2223.94862862958, 
    -2316.69774440581, 
    -2112.16330010733, 
    -1788.82077646629, 
    -1704.78433846092, 
    -1640.12706801873, 
    -1521.49295271204, 
    -1516.17359040913, 
    -2126.28834649884, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3289.06314121088, 
    -3278.51987777659, 
    -3273.10751793873, 
    -3279.59145349244, 
    -3232.09164319353, 
    -3174.18514286738, 
    -3112.6972678805, 
    -3025.55711250262, 
    -2945.94216071425, 
    -2886.36062687001, 
    -2836.05106496437, 
    -2761.04986268115, 
    -1669.07908457789, 
    -168.641907101383, 
    -113.815953263243, 
    -114.284809107209, 
    -161.837352625598, 
    -186.229276520404, 
    -62.2270904537801, 
    -166.088597033348, 
    75.6556345634199, 
    208.709842893337, 
    342.976484369195, 
    821.994138121736, 
    678.175162858966, 
    1645.8340694859, 
    1373.60301307602, 
    1072.60954501674, 
    374.169307100006, 
    131.891482951263, 
    -174.598249048828, 
    -299.312961240896, 
    -226.628083516343, 
    -1562.98968350367, 
    -1870.49228123988, 
    -1936.49002739884, 
    -2244.14641575317, 
    -2328.61494809756, 
    -2386.93768560019, 
    -2534.60893893696, 
    -2678.57767653172, 
    -2757.57811806263, 
    -2798.47808608923, 
    -2781.35889591162, 
    -2860.47015555148, 
    -2866.67087878732, 
    -2859.44156153765, 
    -2878.80595625208, 
    -2886.46375489101, 
    -2906.63431845534, 
    -2927.40739135059, 
    -2948.32031311514, 
    -2939.47364118518, 
    -2953.8965216249, 
    -2962.42036217565, 
    -2925.2365665927, 
    -2868.90652814397, 
    -2706.88775105065, 
    -2580.06137604409, 
    -2383.17708263846, 
    -2342.65013397661, 
    -2219.7433975066, 
    -2157.56634743617, 
    -1885.37244621183, 
    -1660.36640429523, 
    -1745.8544232581, 
    -1572.19077674379, 
    -1434.73868180603, 
    -1296.43016074459, 
    -1655.47130821373, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3266.09913271298, 
    -3273.04282600428, 
    -3271.43497736163, 
    -3219.11312623574, 
    -3197.02079819084, 
    -3139.08954660516, 
    -3052.85465020909, 
    -2994.33437686591, 
    -2920.36770756327, 
    -2850.47585540122, 
    -2789.54594665732, 
    -2048.50315311854, 
    -197.214303060446, 
    -138.201902803888, 
    -49.3151361688621, 
    12.0014780579634, 
    -27.5073298102387, 
    -7.566835472324, 
    32.5193949269024, 
    87.9135907596082, 
    143.45841968874, 
    291.686853156788, 
    154.504549027556, 
    669.569219762234, 
    1379.60212818586, 
    1835.43833161255, 
    1550.97500542003, 
    569.317379659929, 
    705.085037393785, 
    652.55763617128, 
    -108.401093350546, 
    -282.795395401531, 
    -292.346018555187, 
    -1320.8172726519, 
    -1691.9750461557, 
    -2025.33697909604, 
    -2166.50101620459, 
    -2246.76629809543, 
    -2447.65600001558, 
    -2542.45089352598, 
    -2635.07661849788, 
    -2693.28815015086, 
    -2755.87039338354, 
    -2780.59242643247, 
    -2803.21868312105, 
    -2852.76207006098, 
    -2883.39502797228, 
    -2870.95752407642, 
    -2877.71793197171, 
    -2873.99172925789, 
    -2897.07489375919, 
    -2913.79522236891, 
    -2839.5934314621, 
    -2772.315713231, 
    -2892.16524424452, 
    -2850.35410868441, 
    -2720.7189290729, 
    -2659.43434824842, 
    -2457.65624538648, 
    -2419.24592571536, 
    -2378.8633952552, 
    -2248.28300139458, 
    -2307.64564044265, 
    -2045.77117400474, 
    -1719.00203382742, 
    -1758.74781163676, 
    -1588.46982363437, 
    -1388.2643129321, 
    -1464.93358973453, 
    -1132.90168528113, 
    -1075.46042179394, 
    -2296.6467099932, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -3242.48422791416, 
    -3245.72030632814, 
    -3213.88212641837, 
    -3177.34222801695, 
    -3129.92566902186, 
    -3098.80484172825, 
    -3039.51609636501, 
    -2978.29071742076, 
    -2919.86639848562, 
    -2840.24460877763, 
    -2608.79453143454, 
    -381.667659951743, 
    -149.375829344234, 
    -110.079479628688, 
    121.251108013098, 
    122.131409102566, 
    46.4047681011791, 
    80.8067533977932, 
    208.177378123714, 
    86.3973426178078, 
    140.234797991404, 
    395.50048331744, 
    225.271098230883, 
    657.976400736332, 
    1069.28526936667, 
    1857.42185536691, 
    1647.88214810191, 
    637.805238670364, 
    434.371798495039, 
    166.044161350172, 
    -69.2232244094153, 
    -233.877740150868, 
    -511.899087899476, 
    -482.814301335927, 
    -1674.3455553215, 
    -1933.30130215054, 
    -1860.01438134889, 
    -2097.30089956115, 
    -2342.72357570738, 
    -2526.30118816244, 
    -2578.73368334797, 
    -2605.82410484733, 
    -2681.83257612376, 
    -2722.32326252116, 
    -2773.02674361653, 
    -2796.92178348144, 
    -2795.16137527859, 
    -2806.10200208299, 
    -2819.18710405749, 
    -2873.10301944951, 
    -2882.42182708774, 
    -2901.01499554505, 
    -2907.94283647527, 
    -2917.33945149831, 
    -2932.75060515708, 
    -2914.68356500948, 
    -2670.79537799831, 
    -2506.89850010717, 
    -2477.85068599961, 
    -2449.0296644529, 
    -2410.06160754025, 
    -2280.59911101236, 
    -2197.90334751518, 
    -2202.50981579276, 
    -1829.71625873356, 
    -1697.76322267197, 
    -1723.97695760524, 
    -1471.98289404311, 
    -1484.85189834714, 
    -1279.90366015802, 
    -788.036943476249, 
    -1186.5077541048, 
    -2265.19717390139, 
    -2300, 
    -2300, 
    -2300,
  
    -3210.1651497528, 
    -3211.6791563301, 
    -3147.74318463538, 
    -3108.93046660386, 
    -3073.72028770319, 
    -3029.29153753368, 
    -2978.87906451081, 
    -2950.23755658567, 
    -2904.95336357023, 
    -2848.78044615401, 
    -2084.43919485332, 
    -136.387290621391, 
    -168.995820736431, 
    -144.230534341003, 
    175.43584035679, 
    79.0352887063429, 
    450.894134470234, 
    676.956723656403, 
    779.628683903991, 
    699.309698397483, 
    450.599892542586, 
    318.232613989665, 
    279.792180313388, 
    659.819863057756, 
    1444.71062535268, 
    1856.8480463658, 
    1668.95163838727, 
    1373.65711872575, 
    811.478473095172, 
    374.418293603726, 
    199.620131972232, 
    -265.666384352014, 
    -347.766093707962, 
    -237.953792085039, 
    -1255.27440480128, 
    -1876.70159783956, 
    -1937.18311686585, 
    -2057.02501170125, 
    -2268.91015074795, 
    -2474.33677774154, 
    -2447.81932684716, 
    -2487.62453277007, 
    -2549.32396018785, 
    -2615.24644659882, 
    -2693.8731587614, 
    -2739.95089212484, 
    -2750.81119902163, 
    -2755.61558889836, 
    -2783.41594365409, 
    -2819.21153319082, 
    -2869.23205518562, 
    -2876.13003341829, 
    -2890.69998011744, 
    -2910.97330210858, 
    -2862.13000300323, 
    -2753.6088841215, 
    -2705.05668136067, 
    -2618.32253830109, 
    -2532.88975304479, 
    -2535.34757402683, 
    -2350.82384826728, 
    -2242.03446008697, 
    -2192.82176302475, 
    -2249.3106093113, 
    -1936.66695996121, 
    -1699.909531887, 
    -1697.01607334867, 
    -1521.14578014686, 
    -1319.44655695421, 
    -1454.24670076957, 
    -979.128018668622, 
    -936.947398699411, 
    -1303.38525646931, 
    -2113.78560372722, 
    -2300, 
    -2300,
  
    -3126.28193208325, 
    -3141.89720111091, 
    -3103.30195236633, 
    -3054.86575894927, 
    -3037.26268294143, 
    -3003.08592553902, 
    -2953.88107839757, 
    -2905.40878312986, 
    -2845.13281858301, 
    -2668.87000680477, 
    -1405.9677095189, 
    -165.169926958415, 
    -134.399984659835, 
    -88.2688723149809, 
    201.050860606805, 
    582.920104664357, 
    917.006521637201, 
    1224.18562084509, 
    1197.59155924456, 
    1088.48764270471, 
    943.232710920543, 
    539.196423982301, 
    855.20007777027, 
    894.886856002207, 
    1330.72552739706, 
    1659.78759225672, 
    1701.73874767684, 
    1710.70456715207, 
    1009.79057165916, 
    646.039727765276, 
    262.680891914837, 
    -155.266297064069, 
    -287.730834520942, 
    -216.063770518457, 
    -678.13324340702, 
    -1764.41450442393, 
    -1821.03551907769, 
    -2043.28973012756, 
    -2246.13936280937, 
    -2247.92337541912, 
    -2315.2225707461, 
    -2356.91688894718, 
    -2435.67503044239, 
    -2532.49357582767, 
    -2628.51979996189, 
    -2676.12156795147, 
    -2685.78074681879, 
    -2722.00602754634, 
    -2770.59127530806, 
    -2812.14270771364, 
    -2877.77714608631, 
    -2875.1826663642, 
    -2870.95716360675, 
    -2891.52765053197, 
    -2849.57021226701, 
    -2842.38045126647, 
    -2700.45877943221, 
    -2621.19929690644, 
    -2657.70594960177, 
    -2425.46375249882, 
    -2394.59408818808, 
    -2271.98295519787, 
    -2270.079937874, 
    -2146.04854974181, 
    -2106.12098794661, 
    -1780.25637159529, 
    -1705.58929573221, 
    -1607.36577571172, 
    -1439.52296008615, 
    -1457.07770262374, 
    -1161.1857231627, 
    -839.450811448049, 
    -1000.72748374299, 
    -1390.28807741103, 
    -1811.68307302036, 
    -2300,
  
    -3087.99496022531, 
    -3118.42451895685, 
    -3058.91704795983, 
    -3013.42803644093, 
    -2995.94720383801, 
    -2953.02870118418, 
    -2955.31497971555, 
    -2905.28317643493, 
    -2799.50199338223, 
    -1972.86419450478, 
    -259.554384537, 
    -167.559141624682, 
    -89.4595410404654, 
    235.816050945973, 
    370.741224248351, 
    696.824631514765, 
    1181.59262874385, 
    1308.24493162149, 
    1242.13657603846, 
    1125.65397490259, 
    1226.77897006694, 
    1366.83926770935, 
    1043.80726133989, 
    1265.99368118679, 
    1621.67042006678, 
    1496.1430218089, 
    1412.37029142475, 
    1679.00341588413, 
    1229.4892354113, 
    820.076665077333, 
    513.215189678544, 
    35.6547021173009, 
    -154.114133121454, 
    -255.556175477561, 
    -253.642252705268, 
    -1380.15122066554, 
    -1755.08468510029, 
    -1752.11491582002, 
    -1840.07312835318, 
    -1986.2520538706, 
    -2110.5112599611, 
    -2233.75528213826, 
    -2386.43338173314, 
    -2521.39230565395, 
    -2585.66785409549, 
    -2624.03990684244, 
    -2669.66203060342, 
    -2682.92835511553, 
    -2755.38993098995, 
    -2796.40684716031, 
    -2890.20904517094, 
    -2888.69789398638, 
    -2873.3259387043, 
    -2893.47337534393, 
    -2900.18463162105, 
    -2893.42646528118, 
    -2798.06507342126, 
    -2687.22282756536, 
    -2521.6322991007, 
    -2487.85148605227, 
    -2400.69373125886, 
    -2304.9542818315, 
    -2216.20971067969, 
    -2184.05440159848, 
    -2190.38419881139, 
    -1882.634106541, 
    -1677.21256661922, 
    -1745.67126685267, 
    -1565.96776653431, 
    -1476.70781394215, 
    -1394.55630556386, 
    -932.899997288274, 
    -876.830576752498, 
    -1270.55466024606, 
    -1364.35237753805, 
    -1553.60368217307,
  
    -3032.33419529828, 
    -3071.36910303336, 
    -3046.17610426472, 
    -2997.29412346271, 
    -2967.26794214879, 
    -2935.70321409219, 
    -2905.8435014509, 
    -2849.21612859814, 
    -2517.99558740769, 
    -234.985618144911, 
    -180.500662471519, 
    -100.272340906961, 
    -9.62959988627306, 
    323.65933044279, 
    291.209853327158, 
    740.207256782765, 
    1259.36463419027, 
    1328.87726930488, 
    1211.79858003725, 
    1131.77322049371, 
    1192.94885705006, 
    1197.91736273856, 
    1264.00880401372, 
    1097.5902462027, 
    1358.19834875979, 
    1420.18025383516, 
    1045.13590209722, 
    1622.87196553434, 
    1509.55099324977, 
    924.75064936143, 
    599.08869594903, 
    363.885578070085, 
    -99.0701032384381, 
    -236.903548779973, 
    -390.328218897942, 
    -1056.68468882017, 
    -1717.97281131552, 
    -1380.87521980858, 
    -1512.31279796502, 
    -1760.87822450849, 
    -2058.8817909984, 
    -2225.12093214012, 
    -2374.19916338776, 
    -2465.13442569404, 
    -2573.06916267421, 
    -2578.58433766808, 
    -2646.8145297436, 
    -2661.46262960231, 
    -2757.66339432566, 
    -2782.173944249, 
    -2820.04301020333, 
    -2860.54436828682, 
    -2840.47755160444, 
    -2892.42736344802, 
    -2889.07244869629, 
    -2889.58001787585, 
    -2888.97817220827, 
    -2763.33647892216, 
    -2660.80547989763, 
    -2523.53294787775, 
    -2283.56770886874, 
    -2413.9579770557, 
    -2121.43200646002, 
    -2129.66960162839, 
    -2154.02908684025, 
    -2030.96430759066, 
    -1706.34609141248, 
    -1765.11471988212, 
    -1552.19137123851, 
    -1420.5034155082, 
    -1526.06851855852, 
    -1059.0539723361, 
    -794.906067176466, 
    -959.375974298463, 
    -1378.86592066168, 
    -1403.15820840492,
  
    -2985.51461173439, 
    -3024.46190791114, 
    -3028.21126181334, 
    -2958.05372255673, 
    -2927.04462517443, 
    -2898.08268459273, 
    -2857.34432774936, 
    -2769.26681535642, 
    -1004.29786696654, 
    -165.715135736669, 
    -144.137088154091, 
    -84.5084826585837, 
    41.4283992045392, 
    656.424265085116, 
    917.521971391797, 
    868.067115074573, 
    1063.19804249045, 
    1129.26633375623, 
    1051.01858857124, 
    952.333237582867, 
    1230.50485936899, 
    1275.91981554192, 
    1268.55010010654, 
    1311.81976138945, 
    1692.35613982916, 
    1419.96250705356, 
    1148.9565622601, 
    1399.2549892652, 
    1695.36752319337, 
    1237.02587290867, 
    775.192848641283, 
    102.637602353284, 
    -113.61803297767, 
    -258.721430995294, 
    -303.537107145128, 
    -381.154287583896, 
    -1541.30515840366, 
    -1226.91821588087, 
    -1591.38869943651, 
    -1996.2079034957, 
    -2032.62519135854, 
    -2108.65266532941, 
    -2259.38052699654, 
    -2470.87903621456, 
    -2467.89378423573, 
    -2501.90528468082, 
    -2595.92528377589, 
    -2674.45421129592, 
    -2708.82672447213, 
    -2824.48194470037, 
    -2829.04307961117, 
    -2804.56931926048, 
    -2855.95419352533, 
    -2874.46281756052, 
    -2898.94951035862, 
    -2854.57070560605, 
    -2878.83947432669, 
    -2726.10290448743, 
    -2554.64818567017, 
    -2557.17037857927, 
    -2396.44778292016, 
    -2461.40803047684, 
    -2219.06372808476, 
    -2100.05195639889, 
    -2121.21128747818, 
    -2096.74075235365, 
    -1853.16971993954, 
    -1665.76441827413, 
    -1693.18539223666, 
    -1337.22223829929, 
    -1536.67866536618, 
    -1361.79140068302, 
    -944.593863355886, 
    -842.222421626897, 
    -1216.72009183365, 
    -1389.46536453093,
  
    -2951.48445992294, 
    -2974.64422118731, 
    -2989.06705966108, 
    -2973.27965273115, 
    -2926.94639490006, 
    -2871.42815403442, 
    -2802.76521829261, 
    -2508.98106755067, 
    -674.713897337706, 
    -128.658415794373, 
    -150.221050279539, 
    -33.3175065534778, 
    207.172892293897, 
    547.530978989897, 
    742.256469248127, 
    1092.78090053443, 
    1147.53760715668, 
    966.289531814559, 
    778.838126914099, 
    914.756294754558, 
    1118.41703690447, 
    883.930735238856, 
    1008.00681448463, 
    1096.73575826989, 
    1104.69811343613, 
    1001.38431204767, 
    994.64208623837, 
    836.900380432538, 
    1088.18684127483, 
    1191.1671173335, 
    876.604657522372, 
    434.365148048784, 
    -99.6590469836668, 
    -383.031433242169, 
    -426.850482223016, 
    -532.584003401495, 
    -519.346007813804, 
    -1493.50713169828, 
    -1803.25029823841, 
    -1871.39474123349, 
    -1831.90805410832, 
    -2100.72084341017, 
    -2315.67345788151, 
    -2392.18139638185, 
    -2440.90422514332, 
    -2449.86681332647, 
    -2497.63560128719, 
    -2603.2195220298, 
    -2710.63556844577, 
    -2788.93853575225, 
    -2787.72233955751, 
    -2786.9254855063, 
    -2800.03948612363, 
    -2882.65682634821, 
    -2865.47669547189, 
    -2865.38177288607, 
    -2884.97141610174, 
    -2634.89564642313, 
    -2613.79681341805, 
    -2559.45722098526, 
    -2330.32908427034, 
    -2318.64772705215, 
    -2281.77598375275, 
    -2121.52054215759, 
    -2040.12294163549, 
    -2043.50771752984, 
    -1953.71716860507, 
    -1667.63382867042, 
    -1703.12075313555, 
    -1452.55823020465, 
    -1504.11664978574, 
    -1512.63408593395, 
    -929.194951278496, 
    -772.900969134734, 
    -858.938047556438, 
    -1339.1653186247,
  
    -2901.71234787004, 
    -2913.93687837095, 
    -2925.84594788076, 
    -2916.72948986365, 
    -2890.90727201421, 
    -2829.70183967343, 
    -2724.92053752357, 
    -2515.20836066132, 
    -906.35303921074, 
    -148.646805742954, 
    -117.099944655065, 
    16.2124801173323, 
    164.260384582052, 
    436.891331769857, 
    752.315318535847, 
    954.262848489895, 
    1003.19906819548, 
    835.912292540274, 
    710.345123333733, 
    959.977683294795, 
    1254.07901713509, 
    1189.75151437928, 
    1191.64988932337, 
    1170.79978580624, 
    1328.97565428594, 
    1271.54635295462, 
    1193.00175395765, 
    1323.65057678906, 
    1208.14094803181, 
    866.555304190877, 
    566.262191422177, 
    133.698171963749, 
    -110.749507848521, 
    -320.846752773339, 
    -520.118683292778, 
    -503.286102978408, 
    -420.650486564852, 
    -1647.82314632882, 
    -1749.6093870635, 
    -1659.38435777278, 
    -1938.24630204187, 
    -2205.4534248446, 
    -2378.41214245565, 
    -2335.6688686939, 
    -2300.28114963032, 
    -2317.95666404801, 
    -2429.08011718613, 
    -2568.64684604077, 
    -2671.91934771394, 
    -2720.47699060045, 
    -2785.79691228407, 
    -2777.9911396159, 
    -2779.16306772264, 
    -2818.28423645088, 
    -2849.47456105265, 
    -2852.96540031134, 
    -2865.16785535994, 
    -2837.90451839229, 
    -2670.0210049107, 
    -2606.52891784873, 
    -2587.70459811391, 
    -2276.08157830489, 
    -2351.98535730377, 
    -2102.82404405139, 
    -2049.19788774958, 
    -2013.56244875576, 
    -1983.44459663553, 
    -1790.40996540407, 
    -1628.67275555003, 
    -1592.33991050934, 
    -1456.01204212355, 
    -1450.36633442604, 
    -1253.57818222472, 
    -809.245398996658, 
    -860.993907497018, 
    -1025.86116406312,
  
    -2909.91274740768, 
    -2897.65494850902, 
    -2874.28294220483, 
    -2854.91412476543, 
    -2833.31517068109, 
    -2770.21850507337, 
    -2663.5806102176, 
    -2130.20097226338, 
    -1146.03398447583, 
    -317.319558975545, 
    -171.102722258745, 
    10.0697077997317, 
    124.995401170995, 
    589.506799046429, 
    1137.62574393859, 
    1074.95378452826, 
    946.935092212637, 
    666.833727427586, 
    707.169507803067, 
    904.11986231617, 
    1052.65642211846, 
    944.201649323024, 
    814.681404652016, 
    1028.32342191827, 
    1097.1575053387, 
    1145.30726165601, 
    1192.32032656269, 
    1418.15180531809, 
    1503.72333412982, 
    1019.36028493985, 
    534.454366164935, 
    299.687035183627, 
    -101.094833031214, 
    -387.016226197147, 
    -356.756757409416, 
    -205.2822636458, 
    -894.605887708846, 
    -1548.45096590698, 
    -1535.52552009403, 
    -1858.03348745451, 
    -2157.47913233297, 
    -2235.45550687476, 
    -2220.39100833222, 
    -2189.27787010133, 
    -2190.69061689388, 
    -2179.18983587626, 
    -2374.30480895518, 
    -2518.68214189245, 
    -2611.41977841163, 
    -2701.65677143024, 
    -2754.91841909787, 
    -2780.078643047, 
    -2784.4083409838, 
    -2807.12080446523, 
    -2856.50417171534, 
    -2840.18970399795, 
    -2860.30410616235, 
    -2871.8129598483, 
    -2801.55698387086, 
    -2648.11395431126, 
    -2520.53449029698, 
    -2403.73443213929, 
    -2261.25332460478, 
    -2173.38079642608, 
    -2012.88247776352, 
    -1968.81374660718, 
    -1938.44779935796, 
    -1808.41357167277, 
    -1624.30925568755, 
    -1593.56329215841, 
    -1435.67710507383, 
    -1335.81520471861, 
    -1504.52116142862, 
    -857.061581875412, 
    -754.91383208887, 
    -822.701927911261,
  
    -2833.15371926234, 
    -2839.60584921159, 
    -2838.77445592592, 
    -2823.59389431773, 
    -2790.62302432002, 
    -2701.86024264926, 
    -2514.36403359545, 
    -1979.78298364108, 
    -1037.99266844234, 
    -146.669464070746, 
    -112.908148703623, 
    263.57162100951, 
    559.295498462434, 
    876.971128696556, 
    1096.25634924535, 
    1141.70516432947, 
    1136.05038711872, 
    982.903796889077, 
    904.607331356034, 
    927.708890002892, 
    889.515111669047, 
    739.732195650209, 
    735.19045788123, 
    1046.46022310502, 
    985.21767115406, 
    1123.81949052458, 
    1301.79867094068, 
    1179.41229319813, 
    1024.58257764451, 
    569.708726825263, 
    455.974757298107, 
    155.347803256814, 
    161.25885363789, 
    -94.2376758088462, 
    -260.895444419323, 
    -216.562392500719, 
    -1027.8091406913, 
    -1666.39433823401, 
    -1874.01168554975, 
    -1867.10587250132, 
    -1959.07508798836, 
    -2141.56834092092, 
    -2177.74954131362, 
    -2171.0068229513, 
    -2066.93169291156, 
    -2126.42939623313, 
    -2379.51321537577, 
    -2570.96251142786, 
    -2610.24402969548, 
    -2698.38452141603, 
    -2695.03420668513, 
    -2710.5062525494, 
    -2762.7209767238, 
    -2792.96405576084, 
    -2822.38593240121, 
    -2827.21758021646, 
    -2835.14008186913, 
    -2827.28929519226, 
    -2821.66000748962, 
    -2631.03339525246, 
    -2461.70740802077, 
    -2412.38135907044, 
    -2294.82371700411, 
    -2357.15434331776, 
    -2034.70553863969, 
    -1908.43288868459, 
    -1934.3962162099, 
    -1867.09140000979, 
    -1665.89496560433, 
    -1544.75719333149, 
    -1484.77156037846, 
    -1404.69197089354, 
    -1421.45843377706, 
    -1131.85644500492, 
    -752.397718346264, 
    -715.437397408993,
  
    -2783.5683734206, 
    -2795.83514568333, 
    -2813.28292070925, 
    -2790.06919742939, 
    -2749.424138837, 
    -2677.26593547278, 
    -2408.69191489909, 
    -1199.46923064331, 
    -557.456260881929, 
    -186.751425073502, 
    8.70599510955413, 
    287.782998118127, 
    579.281849304747, 
    925.789925860396, 
    1161.54416614631, 
    1320.09466313515, 
    1173.65542351358, 
    1219.93937529321, 
    1264.11448452427, 
    1131.59058341681, 
    909.190524384262, 
    940.720058351455, 
    767.871422155705, 
    830.20316869174, 
    1223.37054163131, 
    1082.55964887903, 
    1356.46977797761, 
    1395.41099509039, 
    880.354420763379, 
    1309.9703311728, 
    1049.10713071065, 
    627.71118449417, 
    765.029263990854, 
    341.685090858483, 
    -197.901298104317, 
    -372.470784160619, 
    -475.745826738279, 
    -1472.60231011232, 
    -1652.14873577259, 
    -1604.90130440946, 
    -1964.57670709454, 
    -1990.71260171615, 
    -2026.24339760912, 
    -2083.82888185644, 
    -1962.41242902356, 
    -2055.14342962695, 
    -2353.38244293999, 
    -2567.08156764254, 
    -2611.77434960992, 
    -2609.91442847172, 
    -2694.76383020416, 
    -2673.06054031355, 
    -2703.02764014301, 
    -2755.56483430425, 
    -2777.72897270519, 
    -2822.43410342431, 
    -2819.83856594175, 
    -2733.98681828583, 
    -2665.07481560275, 
    -2698.49629117447, 
    -2570.99377048402, 
    -2203.47186935442, 
    -2300.5542484638, 
    -2278.55388775491, 
    -2108.32691048241, 
    -1905.5457392369, 
    -1902.33944929407, 
    -1848.66558853269, 
    -1707.02309717603, 
    -1505.57253566968, 
    -1493.51630214507, 
    -1443.55506879886, 
    -1382.71508127791, 
    -1419.16284239492, 
    -823.645058259183, 
    -678.965589286232,
  
    -2699.26372419573, 
    -2732.16434078067, 
    -2698.43544872664, 
    -2743.0002301292, 
    -2670.07967028986, 
    -2619.929357958, 
    -2097.75857849805, 
    -224.444089998457, 
    -248.36912561611, 
    -139.027415478483, 
    6.76400098394883, 
    439.936501762501, 
    919.589621856792, 
    1163.99559062005, 
    1298.18144376441, 
    1426.84467675357, 
    1428.72405190804, 
    1219.23626305729, 
    1291.86750140729, 
    1355.20367558085, 
    1208.0081221526, 
    1144.32491592117, 
    1056.23366644027, 
    686.695010536597, 
    952.960933868992, 
    1119.85740427528, 
    1327.29674050736, 
    1667.82659466136, 
    1359.23510417532, 
    1392.38964073121, 
    1298.58228159325, 
    968.702319103551, 
    281.401601384492, 
    358.765503431622, 
    12.8401642929644, 
    -316.353346082426, 
    -246.137547908411, 
    -768.566515428095, 
    -1489.56497834858, 
    -1623.05950878182, 
    -1959.39464120555, 
    -1835.38158873828, 
    -1815.23004324679, 
    -1912.12840517051, 
    -1837.11706542969, 
    -1972.28902608737, 
    -2367.26229711449, 
    -2474.89280733149, 
    -2502.74620912217, 
    -2583.75716520611, 
    -2589.57408581229, 
    -2640.07461288128, 
    -2684.27084248063, 
    -2726.42472072144, 
    -2777.75337494341, 
    -2777.45820284477, 
    -2802.06836778186, 
    -2815.44929577869, 
    -2654.57961984871, 
    -2737.04688849881, 
    -2562.64342045117, 
    -2520.69178917213, 
    -2386.68602821888, 
    -2143.57526906047, 
    -2021.90111759609, 
    -1930.35363022824, 
    -1845.46322372112, 
    -1855.35252230004, 
    -1648.77824823907, 
    -1449.90122439052, 
    -1468.99025563137, 
    -1398.96222506499, 
    -1390.84434688692, 
    -1394.61200612443, 
    -971.948544885646, 
    -673.918625851895,
  
    -2588.71007207206, 
    -2597.21556776502, 
    -2605.67852677263, 
    -2582.11153860402, 
    -2604.35813960196, 
    -2468.4036629774, 
    -1533.43472661684, 
    -453.444709653951, 
    -123.225367137058, 
    -156.077619329412, 
    21.7659877565385, 
    336.03913659825, 
    965.137833547219, 
    1191.03874920784, 
    1377.46957976714, 
    1498.82029112403, 
    1281.42236640819, 
    1067.51744886956, 
    958.427921478853, 
    1135.63423225087, 
    1332.63873588331, 
    1093.21708901332, 
    939.716419181523, 
    767.777387723678, 
    1199.78852690454, 
    991.441528884187, 
    1436.67270001692, 
    1504.36955040807, 
    1289.63703301612, 
    1304.38851202509, 
    1611.72181787095, 
    886.42103343421, 
    504.839640609892, 
    555.476747066417, 
    253.990205835253, 
    -95.2007822493843, 
    -291.626658664973, 
    -213.857675118783, 
    -450.386391348161, 
    -1055.60129026817, 
    -1674.55534349123, 
    -1593.44805019673, 
    -1643.26826979412, 
    -1679.51911890387, 
    -1733.43231049097, 
    -1888.4764245045, 
    -2231.86755466782, 
    -2279.74064084317, 
    -2334.96632810723, 
    -2446.13369392147, 
    -2549.53653206991, 
    -2590.7608856167, 
    -2662.54788539498, 
    -2714.31826785644, 
    -2769.51409139772, 
    -2800.08616188793, 
    -2810.1555666523, 
    -2816.03302330026, 
    -2801.56484038726, 
    -2746.54633890902, 
    -2555.39585403152, 
    -2311.21900152226, 
    -2343.98710685294, 
    -2115.04743210813, 
    -2067.52483566985, 
    -1967.43507024716, 
    -1775.70393079392, 
    -1816.93370314168, 
    -1740.82113406533, 
    -1358.25447003919, 
    -1376.18860131549, 
    -1412.69506651397, 
    -1398.84124810538, 
    -1367.34878714328, 
    -1251.86049502587, 
    -733.0373696544,
  
    -2496.42788696289, 
    -2457.97684840152, 
    -2452.02574398643, 
    -2397.94052766499, 
    -2511.70435373407, 
    -2126.78755348607, 
    -860.758051219743, 
    -78.9444883246171, 
    -73.3695149170721, 
    -101.246890068054, 
    49.9020026106588, 
    397.447544700221, 
    609.834121302556, 
    1292.95077594958, 
    1425.35326184725, 
    1267.09498194644, 
    1152.58940526059, 
    1020.55450800845, 
    1000.12046291954, 
    1017.50354927465, 
    1397.9767552426, 
    1071.84273408589, 
    1134.32482829847, 
    787.656949495014, 
    855.014795403732, 
    783.442000539679, 
    923.647890191329, 
    917.301354257686, 
    1285.28056335449, 
    1355.17411402652, 
    1591.4663848877, 
    1229.49241316946, 
    1028.34590630782, 
    696.07192310534, 
    202.535348791825, 
    25.9033467895096, 
    -188.765342712403, 
    -357.932291934365, 
    -495.839594991584, 
    -307.596336163972, 
    -681.334279913657, 
    -699.043801558645, 
    -880.497808356035, 
    -1044.34052758468, 
    -1425.27411691766, 
    -1811.67409073679, 
    -2029.2075131065, 
    -2065.16213989258, 
    -2210.41277594315, 
    -2410.10229974044, 
    -2479.66402395148, 
    -2529.14336515728, 
    -2590.04690712377, 
    -2683.46451769377, 
    -2718.25452302632, 
    -2773.77553036338, 
    -2803.9334283126, 
    -2817.87311915347, 
    -2810.53221050062, 
    -2774.66866583573, 
    -2530.09789878444, 
    -2407.28670461554, 
    -2361.53311639083, 
    -2166.35034500925, 
    -2077.46456427323, 
    -2096.44410785876, 
    -1757.39672851562, 
    -1719.04426976254, 
    -1804.68206626491, 
    -1418.54486083984, 
    -1329.72042605752, 
    -1383.06074925473, 
    -1277.3360202187, 
    -1287.08149638929, 
    -1336.52839018169, 
    -937.798812464665,
  
    -2482.88179229702, 
    -2324.78721312793, 
    -2203.45162030911, 
    -2105.84308015112, 
    -2378.91750175929, 
    -1578.51795294784, 
    -165.447251801528, 
    -372.806678434502, 
    -214.522051141617, 
    2.73804636648378, 
    76.7781354267689, 
    673.119032369615, 
    919.539621983236, 
    1097.01994745782, 
    1452.75324274044, 
    1340.9401930652, 
    1080.71124431614, 
    986.9872014899, 
    965.784433627583, 
    1034.17952770135, 
    1094.85007217937, 
    861.457191954267, 
    785.533379378537, 
    652.139885674932, 
    602.457324439174, 
    597.0801585882, 
    771.805799905024, 
    1054.50727120599, 
    1171.04178733014, 
    1240.00001076488, 
    1305.10589698715, 
    1665.86228548159, 
    1177.81556795639, 
    568.441675414698, 
    807.756545563426, 
    455.110945630039, 
    -28.340487254828, 
    -411.165333499035, 
    -522.180859000792, 
    -244.953998300823, 
    -212.203498323447, 
    -258.249339429422, 
    -239.265770308781, 
    -218.229926597365, 
    -325.390748894362, 
    -1462.87094681795, 
    -1664.0684595909, 
    -1767.38660284814, 
    -2077.60260045649, 
    -2275.55225005796, 
    -2354.5989416791, 
    -2402.10331160491, 
    -2468.0395300375, 
    -2601.11428016244, 
    -2689.26035741996, 
    -2714.28489731194, 
    -2779.83578392106, 
    -2810.48310324059, 
    -2778.82269181169, 
    -2782.30338993905, 
    -2568.93267952127, 
    -2398.35619266249, 
    -2304.23711918984, 
    -2229.03224477736, 
    -2108.07125540089, 
    -2054.59072650427, 
    -1788.61349260046, 
    -1689.69593872549, 
    -1748.1271699946, 
    -1526.15427394409, 
    -1224.35623156984, 
    -1322.73197275741, 
    -1324.40433142514, 
    -1308.76414117247, 
    -1258.94710464734, 
    -1169.15826474112,
  
    -1975.96819468602, 
    -1672.55834168096, 
    -1500.27757914202, 
    -1789.10657105654, 
    -2077.8463695052, 
    -1158.78362541583, 
    -95.4441833090274, 
    -103.618768483768, 
    -119.557016609764, 
    137.566150969647, 
    534.697183359112, 
    728.751606342108, 
    652.55910931082, 
    924.898253087367, 
    1322.28934014845, 
    1117.33634796655, 
    968.574382273642, 
    970.920406790089, 
    937.484364047162, 
    896.334431211465, 
    813.33271554603, 
    585.536381985278, 
    488.897971936062, 
    495.342732680471, 
    493.546519865782, 
    652.865896765356, 
    860.118770945379, 
    883.944864048802, 
    962.924160084825, 
    1290.25175170215, 
    1540.541354975, 
    1568.27931724283, 
    1538.3024239193, 
    792.046884536741, 
    314.329874322776, 
    1018.1278465758, 
    105.367062838319, 
    -708.792623598925, 
    -231.714530989677, 
    -266.216598446666, 
    -235.313525224453, 
    -237.189504187692, 
    -231.193490377599, 
    -277.088329259653, 
    -295.713681463432, 
    -358.992463303039, 
    -1170.35723670199, 
    -1690.85929448554, 
    -1958.69406746483, 
    -2104.9112596672, 
    -2215.28466065547, 
    -2288.43499157811, 
    -2382.82202459423, 
    -2511.08039741473, 
    -2605.33175707024, 
    -2691.12161012246, 
    -2711.76438926022, 
    -2732.51118898125, 
    -2730.46319573243, 
    -2793.70925653849, 
    -2627.2543462089, 
    -2466.16698815494, 
    -2202.18182007383, 
    -2148.8682964876, 
    -2069.2315624959, 
    -1867.46223892263, 
    -1773.49900363354, 
    -1670.90040627679, 
    -1652.07795011343, 
    -1591.65581926813, 
    -1205.85306999318, 
    -1300.52316848054, 
    -1206.19920280773, 
    -1187.78068832961, 
    -1124.3236008972, 
    -947.802883562556,
  
    -1644.95593994756, 
    -1464.07648981485, 
    -1267.50389435737, 
    -1524.58395151649, 
    -1784.50241850952, 
    -691.22924095572, 
    -34.0223712200277, 
    -90.6512095717275, 
    -100.70859622635, 
    121.603477995447, 
    415.636118714782, 
    839.356941505082, 
    849.168063976465, 
    929.032407822562, 
    1148.21918654148, 
    995.991046986681, 
    1129.24625662433, 
    970.357581571128, 
    835.284022315218, 
    759.101379796078, 
    674.121508189305, 
    540.97456335087, 
    479.12592803938, 
    524.31078355283, 
    607.835073054571, 
    764.033859295648, 
    920.350990611522, 
    974.08015536728, 
    731.815738109831, 
    1169.50143536849, 
    1281.60734703346, 
    1299.61335798821, 
    1205.9247704791, 
    979.630153549215, 
    905.6289411846, 
    820.942497287587, 
    2.82838661913518, 
    -698.550527690101, 
    -251.222885027178, 
    -292.20879066698, 
    -274.568453426724, 
    -274.462056598898, 
    -288.602411872463, 
    -351.922525638696, 
    -389.176891745539, 
    -379.617001681952, 
    -340.90582141684, 
    -938.118480438888, 
    -1766.46524724501, 
    -1926.67734808671, 
    -2029.30058961806, 
    -2127.21836683865, 
    -2275.10646140856, 
    -2408.49740193913, 
    -2488.2969671337, 
    -2584.66426939073, 
    -2653.80099118223, 
    -2723.04651124961, 
    -2722.0013967687, 
    -2715.04873264223, 
    -2683.01011488552, 
    -2465.32307203406, 
    -2262.06295407286, 
    -2166.90811509221, 
    -1990.59932123507, 
    -1905.17846435342, 
    -1734.52752847874, 
    -1590.14427873669, 
    -1566.32038423169, 
    -1573.48112253699, 
    -1228.61430534884, 
    -1209.73469996265, 
    -1141.21061248608, 
    -987.221525220026, 
    -805.96066014203, 
    -589.924862168536,
  
    -1364.07488261839, 
    -1169.27454722235, 
    -1081.80992934685, 
    -1375.31722829377, 
    -1643.3654540298, 
    -252.520720818276, 
    -218.161409893872, 
    -298.717433527897, 
    -39.5466698004813, 
    158.420908664136, 
    429.974573923512, 
    1150.80024884983, 
    1253.92359447586, 
    1040.56269467344, 
    1001.54107279847, 
    680.161849855975, 
    853.50132557526, 
    807.010811245053, 
    704.815229956272, 
    659.240974844903, 
    623.33003147719, 
    585.570096749608, 
    538.122212126968, 
    550.501537421249, 
    582.212124729475, 
    594.18870913515, 
    720.130590603305, 
    569.340001498195, 
    648.409964054189, 
    1034.77352330292, 
    1144.67834230019, 
    1073.55340475358, 
    869.699170171346, 
    895.663670530242, 
    482.615674577387, 
    126.555615111136, 
    26.9008742736365, 
    -467.561246767285, 
    -267.49432086197, 
    -375.248505386233, 
    -349.683175218332, 
    -369.668255330734, 
    -452.578629142361, 
    -435.640254589906, 
    -463.111743961177, 
    -426.632899541737, 
    -391.628777199603, 
    -402.631621665143, 
    -1281.35854953881, 
    -1643.3347477758, 
    -1774.56390360355, 
    -1916.92008907237, 
    -2099.78825260517, 
    -2249.01144805601, 
    -2324.69474131209, 
    -2400.10892608745, 
    -2530.09065743817, 
    -2644.49756549694, 
    -2703.7394671296, 
    -2685.3555444459, 
    -2688.86352716768, 
    -2503.50647437425, 
    -2256.83951417383, 
    -2179.51517577988, 
    -1910.93656019187, 
    -1811.82184868243, 
    -1617.74639210802, 
    -1509.69998888313, 
    -1464.17202162449, 
    -1458.97273543167, 
    -1197.81618104189, 
    -1112.65728522255, 
    -952.230674162689, 
    -637.597749118438, 
    -366.546567833568, 
    -303.993953807357,
  
    -1148.61492499579, 
    -1100.04205240248, 
    -1039.10675819457, 
    -1381.2365178261, 
    -1305.83126328694, 
    -133.664718254146, 
    -186.756396115291, 
    -83.941207588319, 
    -9.64202815074022, 
    223.669974550286, 
    871.270385588408, 
    1151.21394777886, 
    889.805892209592, 
    935.286896059521, 
    827.512050188668, 
    585.571287481942, 
    747.180902658358, 
    548.397098203788, 
    458.951742755338, 
    458.429874445796, 
    580.782864313242, 
    641.98827432972, 
    608.483342639543, 
    594.418141936402, 
    562.345795301415, 
    450.048649133254, 
    647.541146640415, 
    839.324226302504, 
    913.191209346692, 
    1078.94142942012, 
    1470.67814658444, 
    1441.60660970758, 
    968.488773811569, 
    698.435146165188, 
    141.730678560489, 
    365.865311973976, 
    30.6731653157437, 
    -25.5337187119856, 
    -215.126923098676, 
    -321.046523103789, 
    -443.72364230439, 
    -505.008752517445, 
    -732.625353959482, 
    -779.720694290966, 
    -591.699704656141, 
    -456.263028891329, 
    -392.222251806654, 
    -331.95894005958, 
    -332.536619098827, 
    -1006.70756288125, 
    -1607.83675026546, 
    -1803.21814169889, 
    -1947.44286788137, 
    -2014.74458157495, 
    -2159.03223179116, 
    -2299.13690739169, 
    -2446.28580374894, 
    -2554.87642831151, 
    -2616.23856882606, 
    -2698.71691412675, 
    -2676.19539612431, 
    -2536.21644809291, 
    -2329.05216366553, 
    -2119.35736398387, 
    -1891.6480412841, 
    -1678.19931226775, 
    -1481.73031486349, 
    -1418.79144905663, 
    -1315.13580670843, 
    -1281.02408344401, 
    -1153.57896982088, 
    -949.414801807979, 
    -634.646633536922, 
    -385.256098252793, 
    -326.817221728044, 
    -320.488669533212,
  
    -1097.68593036101, 
    -1077.68111941689, 
    -1109.56653771822, 
    -1424.19622419983, 
    -982.869622643824, 
    -70.5284259316634, 
    -86.0157566545783, 
    -109.644206021428, 
    -0.631521467832885, 
    398.231326975722, 
    768.496167549237, 
    568.424160383848, 
    486.870255281246, 
    536.319385840405, 
    705.396867228782, 
    481.746514127077, 
    715.495003131039, 
    460.304938172172, 
    537.577505139462, 
    530.552082561567, 
    503.278541052329, 
    589.934036280514, 
    678.47398083421, 
    702.999114383643, 
    709.651056877045, 
    780.152132980503, 
    784.785178138588, 
    758.615466306885, 
    777.866834437592, 
    1007.64112787364, 
    1165.36819562239, 
    1084.89876273605, 
    879.744881863824, 
    978.261010045035, 
    1218.86104128369, 
    1004.09459246286, 
    353.132994022774, 
    181.520782721133, 
    -203.026550559955, 
    -311.954269127243, 
    -567.863402858963, 
    -490.008605704996, 
    -645.156699877971, 
    -732.91488335621, 
    -454.551052102047, 
    -290.831412764974, 
    -311.125710763964, 
    -349.574976576137, 
    -391.105274640434, 
    -382.655001568768, 
    -1021.5696041026, 
    -1620.11499031981, 
    -1681.26426655768, 
    -1811.67450122043, 
    -1963.45607819936, 
    -2080.06316233055, 
    -2311.18924667854, 
    -2445.00299581461, 
    -2547.17711623172, 
    -2615.90740508862, 
    -2590.43081753892, 
    -2540.22951696381, 
    -2309.74458037886, 
    -2094.84429422445, 
    -1847.52144076869, 
    -1591.32809359389, 
    -1475.93747207966, 
    -1338.48053921724, 
    -1179.53240783965, 
    -1108.65212245484, 
    -975.024023382817, 
    -598.039162006781, 
    -294.080593442328, 
    -269.572615334061, 
    -327.725820060807, 
    -397.875226122267,
  
    -1133.7382379, 
    -1141.25494664994, 
    -1175.84090325333, 
    -1160.1446891178, 
    -599.955669620932, 
    -55.7722079793923, 
    -64.7302838909664, 
    -74.1440887056037, 
    -12.1134328468388, 
    363.117831656277, 
    384.528860132746, 
    471.490293496391, 
    368.380367210696, 
    599.350097844207, 
    564.055521231348, 
    876.187953560246, 
    868.358859815098, 
    668.214998473781, 
    735.260910649317, 
    699.085904897796, 
    537.674549397537, 
    609.941260471323, 
    738.321702211729, 
    809.693311240613, 
    718.985722694523, 
    781.633312272331, 
    765.880272851414, 
    747.361606533828, 
    1044.69792646043, 
    1053.76239732185, 
    1049.3909640937, 
    1036.56971737306, 
    1018.29346583965, 
    936.75645287867, 
    1154.73737291633, 
    1098.05545782108, 
    487.766672456911, 
    -35.4690333357861, 
    -205.614462823644, 
    -283.23974662345, 
    -464.084524742033, 
    -701.611946046152, 
    -605.76748994697, 
    -437.666020067648, 
    -414.921351771338, 
    -496.053340834974, 
    -549.264429978805, 
    -591.130638284887, 
    -563.046570328288, 
    -398.823859578951, 
    -832.17184773752, 
    -1342.1909205489, 
    -1407.82425816996, 
    -1534.59143811404, 
    -1741.12312439922, 
    -1937.78038211152, 
    -2152.38904625358, 
    -2348.66880680439, 
    -2458.51045867817, 
    -2497.61973214657, 
    -2507.35534049415, 
    -2479.28967268069, 
    -2246.68963930615, 
    -2002.94635293411, 
    -1693.66918453203, 
    -1506.22489891607, 
    -1402.04953489912, 
    -1264.06360218693, 
    -1027.90012951687, 
    -908.404484107004, 
    -662.84407700456, 
    -348.035132473286, 
    -333.97371692807, 
    -227.675045032651, 
    -210.356281842256, 
    -293.074143818751,
  
    -1179.30975704044, 
    -1134.51708171029, 
    -1053.62312156276, 
    -835.708310023663, 
    -269.418619756069, 
    -153.768459754723, 
    -92.8962159066024, 
    -49.0095148305474, 
    35.3157918818997, 
    128.14834566319, 
    166.036044734858, 
    765.327902175543, 
    312.318218380705, 
    294.843525272461, 
    630.751378186472, 
    1071.19102119198, 
    1018.60248132516, 
    827.348572759853, 
    836.904603460469, 
    734.783005469856, 
    668.885698427411, 
    595.445082293912, 
    648.877573498151, 
    745.75793697105, 
    770.936076011531, 
    920.432002154071, 
    980.266034347348, 
    828.026244946315, 
    881.564977929945, 
    889.268068328547, 
    1094.21530332491, 
    961.781409909715, 
    772.562128961959, 
    1055.68705930635, 
    939.76558676759, 
    450.866038729325, 
    257.898018946971, 
    -18.117408533246, 
    -71.4977209864371, 
    -210.50795689035, 
    -304.234193769842, 
    -670.331624209416, 
    -555.351918766238, 
    -393.267412209163, 
    -333.801384792349, 
    -409.433395714668, 
    -567.410767686593, 
    -494.731849751571, 
    -309.579893883235, 
    -318.995653530517, 
    -888.299431342693, 
    -1084.94972850974, 
    -1078.82660019758, 
    -1316.17587387922, 
    -1605.95797358702, 
    -1851.13671324795, 
    -2106.95100107225, 
    -2262.51122520592, 
    -2367.28569869739, 
    -2434.9967080316, 
    -2403.34314245072, 
    -2381.91909718273, 
    -2297.97084597324, 
    -1997.54709644894, 
    -1595.57246781677, 
    -1399.45046819364, 
    -1293.6949995325, 
    -1119.69789034682, 
    -898.854145208103, 
    -734.406547529297, 
    -436.899037992296, 
    -339.561952482012, 
    -338.241792975722, 
    -314.976429763059, 
    -260.26472210003, 
    -203.298243549342,
  
    -1159.88608632189, 
    -1037.36247983038, 
    -884.798171492999, 
    -492.214799028757, 
    -283.272827584158, 
    -411.871353820084, 
    -293.798524096194, 
    -51.9665710133107, 
    68.1450618400016, 
    72.935563970121, 
    201.204184405077, 
    74.9500553327605, 
    583.591959095743, 
    670.915551880836, 
    720.864541441436, 
    1012.01865386108, 
    876.599389190501, 
    739.317483703336, 
    851.703493261391, 
    752.97949511794, 
    590.173641952394, 
    480.329392162975, 
    492.472280363487, 
    571.498888773987, 
    653.794975203866, 
    817.827299000565, 
    717.811816549776, 
    753.355721083895, 
    872.481964111327, 
    628.529877281401, 
    836.189994282311, 
    952.929932956332, 
    939.239343846099, 
    1063.54323223323, 
    574.167731734698, 
    314.167903524228, 
    25.6061079070956, 
    186.42336362634, 
    0.0134878037426707, 
    -127.162555980789, 
    -240.010619337588, 
    -318.05385686996, 
    -735.248900640985, 
    -514.077608593367, 
    -231.558884329116, 
    -247.466425529386, 
    -348.916031050388, 
    -198.108421690919, 
    -212.377595173151, 
    -320.161674772905, 
    -508.431359747082, 
    -633.540365332312, 
    -886.548579798033, 
    -1146.14534551913, 
    -1532.68934304984, 
    -1718.16876102802, 
    -1975.17815535012, 
    -2146.5100719627, 
    -2267.0062819734, 
    -2275.26633223547, 
    -2268.01920495455, 
    -2301.219535016, 
    -2234.33716995906, 
    -1906.14681024327, 
    -1285.46171089675, 
    -1299.51513905968, 
    -1200.78220481061, 
    -1013.48781803554, 
    -811.563195197604, 
    -652.574063274385, 
    -371.983082415672, 
    -313.124787086068, 
    -307.006218272654, 
    -323.432362128212, 
    -252.00891497314, 
    -218.935219966551,
  
    -1090.06584570736, 
    -921.35462538152, 
    -365.134780260103, 
    -175.825712955811, 
    -88.1462480517278, 
    -114.571755123028, 
    -466.369548126938, 
    -97.2975114243571, 
    48.9926916535726, 
    242.806607429019, 
    60.2974397775742, 
    175.165183385574, 
    106.201597954893, 
    421.487898793487, 
    906.571237758454, 
    898.735446438677, 
    737.25577293131, 
    648.498770437209, 
    919.642096652964, 
    836.13346398878, 
    568.250183250709, 
    464.597384274474, 
    437.558034646952, 
    569.055516335891, 
    681.44007649694, 
    659.493085769363, 
    580.926827826935, 
    897.324093740704, 
    680.693167503842, 
    490.58173201199, 
    827.328981252164, 
    891.061182848682, 
    834.997833063989, 
    582.426001109845, 
    584.789411017236, 
    442.038318804909, 
    419.31409856321, 
    656.762417416293, 
    197.935190640803, 
    -21.29338841509, 
    -141.199086388975, 
    -225.815821353959, 
    -328.899710741714, 
    -300.626705148315, 
    -195.627032560837, 
    -193.984519422388, 
    -218.645523167403, 
    -215.679760263321, 
    -218.246542216149, 
    -241.130846474232, 
    -284.815206863044, 
    -311.036285930091, 
    -465.384682440676, 
    -895.424204323352, 
    -1332.18570879245, 
    -1607.37771418487, 
    -1791.02076316227, 
    -1911.08657455871, 
    -1954.46887642752, 
    -1981.35772949423, 
    -2082.07156983789, 
    -2180.90363703917, 
    -2068.6938018628, 
    -1908.62557621152, 
    -1459.37813944886, 
    -1199.48155145763, 
    -1165.26255181495, 
    -954.636535294245, 
    -715.148747007361, 
    -428.81082105049, 
    -305.060583646461, 
    -280.071237925051, 
    -275.589338663578, 
    -281.689445346093, 
    -269.861780023521, 
    -213.974574504481,
  
    -974.734789276976, 
    -518.461007787821, 
    -254.164385768895, 
    -140.637915317583, 
    -144.01590671518, 
    -188.03018397153, 
    -459.554752371215, 
    -189.249977338219, 
    -0.605989593676771, 
    259.651408743349, 
    263.028109536596, 
    343.669251765545, 
    339.280911124171, 
    829.313548644476, 
    988.823208030369, 
    1001.69461308188, 
    733.605193664619, 
    569.66410482477, 
    677.459021368588, 
    822.280000462374, 
    649.130762892633, 
    567.761484357571, 
    470.686634794195, 
    457.667837068187, 
    456.28800413296, 
    515.428265587612, 
    597.407542605682, 
    595.799800911246, 
    434.300971660207, 
    676.901120817008, 
    778.228786045597, 
    476.382985024274, 
    409.726220330631, 
    530.042913618439, 
    561.115205267105, 
    528.416696042253, 
    657.72418963869, 
    855.798958021208, 
    341.708092432136, 
    13.7715911566189, 
    -41.5234240951619, 
    -114.935766310867, 
    -212.49902342682, 
    -375.211803496085, 
    -212.773422700425, 
    -186.785073700036, 
    -202.868531569923, 
    -213.14384131736, 
    -306.466965264197, 
    -263.744808771575, 
    -269.022315558234, 
    -246.517031145255, 
    -241.913924457512, 
    -376.439583973814, 
    -944.876190638352, 
    -1328.07487511715, 
    -1530.29482459808, 
    -1516.66187384627, 
    -1467.34158877108, 
    -1459.79806691134, 
    -1612.83165410331, 
    -1704.78731296791, 
    -1821.92639647138, 
    -1801.84131214787, 
    -1543.38885380146, 
    -1270.28897969586, 
    -1043.26060583236, 
    -878.883741269853, 
    -517.617773963778, 
    -318.801729020717, 
    -229.050519475477, 
    -210.106212045684, 
    -214.409482891855, 
    -206.423804115474, 
    -217.182505352366, 
    -259.081398153359,
  
    -845.501920300661, 
    -305.792799288588, 
    -264.717475933831, 
    -148.384103661822, 
    -129.603791298818, 
    -128.069781679321, 
    -351.21351183969, 
    -106.433502052025, 
    38.2960580153523, 
    131.797843364962, 
    155.448583058256, 
    432.628729137833, 
    490.032887995984, 
    880.906156319918, 
    921.521328275709, 
    916.294498601657, 
    684.609291102289, 
    562.379071507982, 
    537.553335960874, 
    599.436321365337, 
    701.975617523022, 
    655.33286548542, 
    699.571538987115, 
    515.438719020046, 
    428.031101730875, 
    452.14969102319, 
    351.31668875118, 
    348.408777879842, 
    339.35022849225, 
    372.203717128154, 
    467.362746154338, 
    573.085793455666, 
    485.722931566051, 
    430.044503475756, 
    357.668574291539, 
    335.568660825793, 
    541.095561028595, 
    589.578029081504, 
    106.370182890642, 
    9.75171972349139, 
    27.6087513756594, 
    20.5112075600102, 
    -107.268926745432, 
    -53.4764308276561, 
    -278.061721932044, 
    -44.6596378760117, 
    -188.338239349415, 
    -255.976417947321, 
    -269.511523085505, 
    -304.448270274438, 
    -325.185558135405, 
    -272.115612841668, 
    -219.61259347247, 
    -256.760312912313, 
    -340.446753977124, 
    -605.950302094111, 
    -1086.58061701827, 
    -1102.37341204362, 
    -1063.33966577066, 
    -982.467391267196, 
    -1081.768309983, 
    -1232.10439851596, 
    -1476.96167197232, 
    -1564.76951170234, 
    -1491.40685085113, 
    -1222.67663152167, 
    -995.969480311617, 
    -689.550690790839, 
    -378.023857654942, 
    -266.282363084235, 
    -195.776979354567, 
    -180.301096050096, 
    -188.085760573657, 
    -175.178992618505, 
    -179.644638838987, 
    -247.190341022487,
  
    -829.431029171319, 
    -428.499902838427, 
    -273.982618987627, 
    -155.481610999796, 
    -106.573275923863, 
    -75.3903801096779, 
    -259.963228304734, 
    -117.605540490233, 
    48.4273283466924, 
    375.88434454735, 
    452.612276147758, 
    364.225907358847, 
    464.718811124869, 
    618.377664384489, 
    829.904767556526, 
    757.045277235621, 
    625.701728598668, 
    532.33800292576, 
    603.794443692233, 
    635.010099609646, 
    718.975014698333, 
    734.108261125486, 
    693.418518869499, 
    483.373797037566, 
    334.010275829013, 
    396.829139119966, 
    343.041717849683, 
    425.656408282167, 
    386.158875242192, 
    326.86885342486, 
    403.684035468875, 
    539.175315540818, 
    460.153040703308, 
    404.373816905603, 
    338.26710414566, 
    343.630882425511, 
    431.7730210316, 
    414.822187968356, 
    355.830768828697, 
    643.340013027733, 
    615.928581203633, 
    579.382510006907, 
    333.157664953662, 
    411.898899573895, 
    131.94855568417, 
    108.307644983422, 
    -65.2622934290147, 
    -156.513083194164, 
    -241.470573937906, 
    -280.668784441633, 
    -267.471123258583, 
    -333.275499119602, 
    -269.268710301946, 
    -292.053498403757, 
    -258.721336947845, 
    -299.631528796701, 
    -419.284146371906, 
    -488.257308541316, 
    -423.315558024503, 
    -422.166346358822, 
    -470.762171225208, 
    -562.814126111889, 
    -1014.02393793018, 
    -1291.02133544375, 
    -1378.72372316913, 
    -1203.55802490302, 
    -995.305914858554, 
    -674.607877938505, 
    -368.36115080779, 
    -227.636339258105, 
    -169.901932298802, 
    -160.345276929763, 
    -155.880021878079, 
    -142.237539754869, 
    -139.818545833814, 
    -162.938509256548,
  
    -850.555126801049, 
    -694.45713091057, 
    -437.925656851571, 
    -142.94831109127, 
    -90.288035660815, 
    -72.9484233023202, 
    -191.333491623335, 
    -188.091557177025, 
    27.2211599312601, 
    449.511996817078, 
    562.114457569357, 
    659.933612631256, 
    578.724380228314, 
    629.313571430133, 
    818.996601553271, 
    695.249937324482, 
    622.242797603799, 
    576.931659976152, 
    557.788749532496, 
    536.631467453976, 
    644.723996503085, 
    716.849493507306, 
    620.530230215654, 
    470.309368445385, 
    367.93227007568, 
    374.945848424384, 
    451.880499264161, 
    556.844043078109, 
    559.056717568258, 
    523.146614356647, 
    590.86153477651, 
    582.581973136741, 
    435.095096635123, 
    366.247705675317, 
    313.461648174257, 
    289.156839876932, 
    371.005063367717, 
    519.654538110817, 
    533.700214800348, 
    785.033556785456, 
    1027.85315804306, 
    1049.78883471174, 
    174.778889486271, 
    198.438991002246, 
    545.863901823924, 
    283.908830324458, 
    163.631901764529, 
    2.66889519387123, 
    -179.229459578886, 
    -280.334033385104, 
    -278.596588690096, 
    -264.323240521507, 
    -294.342385209822, 
    -300.688437706412, 
    -282.978456012346, 
    -312.008379411857, 
    -294.638929023188, 
    -299.312834616872, 
    -328.175921052461, 
    -398.273995902477, 
    -408.081385276085, 
    -387.919063098219, 
    -406.041450504758, 
    -969.569383106465, 
    -1172.96066041542, 
    -1046.65013006366, 
    -914.674593499365, 
    -708.058479949848, 
    -418.632232845428, 
    -203.375668419968, 
    -163.666149564446, 
    -144.341486239887, 
    -134.965714658628, 
    -110.912700083862, 
    -98.9271470814236, 
    -86.2990972704738,
  
    -814.163299654525, 
    -734.727817291909, 
    -517.496894229833, 
    -126.425668230516, 
    -134.566871557632, 
    -112.383113281191, 
    -131.559857290509, 
    -79.6763694214222, 
    28.8069615946094, 
    504.666570460532, 
    593.538554303724, 
    520.350425959429, 
    498.953717726206, 
    576.393248460859, 
    706.371678265852, 
    668.560410229381, 
    593.251402390364, 
    529.327653797315, 
    480.432428857647, 
    400.006480564061, 
    522.775592628811, 
    519.512977266897, 
    553.918917152942, 
    465.282966348918, 
    376.19905455569, 
    351.640827097791, 
    469.113135667824, 
    518.89713135278, 
    480.010023806955, 
    563.884391964082, 
    624.303404779205, 
    516.221838149085, 
    302.977288309161, 
    351.499637633663, 
    303.896960229648, 
    218.40891138143, 
    256.784478763185, 
    509.871619528914, 
    495.253749766249, 
    653.670659525527, 
    876.686711361531, 
    1010.44873140854, 
    654.330414997364, 
    75.8243742824722, 
    878.289997686066, 
    766.567639366921, 
    305.198902888375, 
    571.059203533415, 
    -54.1768880133387, 
    -309.901525345789, 
    -256.610839801031, 
    -272.560685250687, 
    -301.946149588966, 
    -300.070343602812, 
    -294.68907981864, 
    -282.405856325805, 
    -260.171646404374, 
    -318.387875709662, 
    -386.779300839211, 
    -422.65380073368, 
    -422.805924081322, 
    -377.806316802908, 
    -319.957617602717, 
    -637.909327610604, 
    -915.494162966392, 
    -973.902167710049, 
    -799.911714107431, 
    -643.391260290198, 
    -419.949312220762, 
    -217.912832371197, 
    -167.841416364287, 
    -131.467035842502, 
    -109.159769169293, 
    -89.0579012713796, 
    -72.0390926117588, 
    -80.0348703078964,
  
    -776.480781862743, 
    -716.615330789017, 
    -378.529269505719, 
    -106.451243827751, 
    -105.809439486111, 
    -100.860984778751, 
    -123.47126519373, 
    146.665092720301, 
    398.915709693122, 
    770.58155838988, 
    435.405634342891, 
    611.581271223894, 
    448.310019767549, 
    380.766043044689, 
    743.169859754815, 
    653.643069926195, 
    508.718556928473, 
    603.931887260345, 
    473.048671478921, 
    428.803967363758, 
    428.453022507243, 
    489.290655843087, 
    430.220626292808, 
    406.869189318988, 
    368.780440946709, 
    226.646926061835, 
    335.492389362841, 
    308.687058221317, 
    367.985963537336, 
    456.22645335181, 
    342.959587366287, 
    412.746238238597, 
    282.536452815623, 
    381.595624285077, 
    158.983031098811, 
    196.568459603717, 
    289.839350530575, 
    388.555554269273, 
    476.296980722221, 
    508.460715200972, 
    684.128779087728, 
    916.938021977026, 
    776.804787263088, 
    60.0826600540409, 
    539.250633882633, 
    1073.14510731628, 
    1164.82272762627, 
    899.82653143051, 
    158.437697031461, 
    -207.91647781209, 
    -177.439547539824, 
    -269.322259695773, 
    -310.13593887295, 
    -306.327679607396, 
    -299.856418720685, 
    -289.470768081648, 
    -275.558236586687, 
    -311.952406862949, 
    -414.630729448889, 
    -465.470199495255, 
    -442.166590674593, 
    -321.889942053849, 
    -297.926726825026, 
    -344.599638833177, 
    -513.679726962677, 
    -621.949912059478, 
    -718.899705115782, 
    -608.410341004374, 
    -435.527009697002, 
    -240.551975876058, 
    -176.267573099253, 
    -123.929747607113, 
    -96.0372854587344, 
    -72.5552489375744, 
    -29.0224495556143, 
    -30.5412121235577,
  
    -740.247630940572, 
    -677.615130314501, 
    -325.513174326127, 
    -104.291587418431, 
    -115.430317991926, 
    -95.7971911360935, 
    -169.848924256654, 
    238.631696508816, 
    416.959230254253, 
    1210.4434583948, 
    1003.91905408906, 
    713.134972900192, 
    1220.86285084281, 
    1189.52863949972, 
    921.563283409811, 
    753.789648323019, 
    566.744716221383, 
    617.16067519407, 
    506.24812940574, 
    512.916979551584, 
    478.19563480561, 
    416.732930259233, 
    361.027920111029, 
    344.16543412075, 
    267.593409236039, 
    229.417100175898, 
    205.640742386307, 
    225.135369408704, 
    241.262965344367, 
    254.203667498647, 
    206.085538014051, 
    290.117390627286, 
    237.936602909645, 
    298.979504998557, 
    182.34370211124, 
    251.13349646283, 
    347.868414657781, 
    181.527475130649, 
    495.320136477136, 
    413.789438066129, 
    385.446550136447, 
    170.693213719145, 
    540.090652841759, 
    982.711081364939, 
    1172.44828271814, 
    1011.06836402271, 
    1301.37082223582, 
    902.207241951131, 
    719.063548076341, 
    519.673045291894, 
    44.5227475323916, 
    -248.709233737872, 
    -325.914765224475, 
    -308.420781284003, 
    -300.412164741508, 
    -298.560266949695, 
    -298.277831740769, 
    -309.908000565857, 
    -433.491377583811, 
    -491.503695185748, 
    -432.949676193287, 
    -296.939844223313, 
    -297.444446106641, 
    -307.974505780125, 
    -378.219611784111, 
    -470.657896928264, 
    -541.018614911015, 
    -620.332433224258, 
    -451.803361510376, 
    -265.400271568427, 
    -236.978110179924, 
    -200.208371189113, 
    -124.15276471124, 
    -66.1614771994604, 
    -33.8336928451446, 
    -6.39979241630749,
  
    -705.046541314376, 
    -617.090352399084, 
    -194.16306791487, 
    -122.081994127186, 
    -117.654790993633, 
    -75.0474929852279, 
    -120.925751669007, 
    124.371804746782, 
    331.753064882856, 
    852.227871346974, 
    618.598065118888, 
    1202.00683706524, 
    1523.85923608179, 
    1106.43604766401, 
    1223.58485716748, 
    883.817273642954, 
    726.452316224377, 
    724.230891203159, 
    610.347495725148, 
    615.260160080932, 
    484.297162477809, 
    380.39995372469, 
    337.787802466619, 
    360.528985048062, 
    213.336151022659, 
    179.760859302549, 
    129.906525616148, 
    163.319909517601, 
    224.026050161808, 
    153.031528660858, 
    147.584558798779, 
    149.551150241864, 
    232.495852603893, 
    165.888404886773, 
    237.858970763838, 
    378.868322203705, 
    247.375205085898, 
    178.887036501893, 
    364.438225100049, 
    355.167429694402, 
    349.28322008823, 
    509.10098631839, 
    1151.03431852027, 
    1488.28396850791, 
    1868.4148208943, 
    1439.19487517252, 
    1287.34929683469, 
    1403.27773593337, 
    1493.49164501844, 
    986.435403163866, 
    353.509507472948, 
    -124.928711372151, 
    -218.356995186373, 
    -284.60718642317, 
    -327.852670727224, 
    -309.05610804969, 
    -301.020554391961, 
    -304.960937717861, 
    -436.458322352018, 
    -451.082529800602, 
    -414.551626839802, 
    -325.787860379107, 
    -301.102555551561, 
    -298.393563901724, 
    -314.037921610766, 
    -441.965294392618, 
    -487.825773036226, 
    -561.45322392582, 
    -578.77862968317, 
    -327.864836087289, 
    -203.482266198612, 
    -156.481628635829, 
    -127.619176434242, 
    -75.1855984940912, 
    -45.216385427541, 
    -14.5198249058665,
  
    -648.12153423006, 
    -509.148155421721, 
    -122.340397582743, 
    -110.425415551676, 
    -100.771452911223, 
    -89.4667140772734, 
    -58.8121481261246, 
    353.064898761094, 
    920.235107447502, 
    1253.26791933749, 
    1524.12535344687, 
    1453.02756494263, 
    916.652958621102, 
    1261.45249539126, 
    1012.6479926371, 
    966.437671229926, 
    840.854498962539, 
    698.134906063955, 
    742.093262333885, 
    648.344959869897, 
    542.494711736015, 
    370.866355767843, 
    303.552293138835, 
    329.063818210718, 
    363.68949357446, 
    201.575743432808, 
    134.310907061663, 
    129.620929632582, 
    117.616835918833, 
    155.007896782169, 
    92.6263327069938, 
    157.978764509433, 
    243.149012404352, 
    131.105429101498, 
    275.297799728752, 
    301.701678661591, 
    218.097297726126, 
    150.767948684607, 
    223.201535672384, 
    339.089555097454, 
    437.031903129143, 
    672.32793129198, 
    1181.32713561363, 
    1755.09726779164, 
    1964.75813655704, 
    1791.60080299505, 
    1732.43937269597, 
    1829.0828574972, 
    1535.05753243544, 
    1309.5721131738, 
    996.11013483814, 
    277.571225842054, 
    -166.868812616569, 
    -270.035381492282, 
    -314.940118321913, 
    -333.391411019866, 
    -302.38755181068, 
    -361.077266167687, 
    -468.404183514842, 
    -454.647222576589, 
    -378.351000355445, 
    -309.226989323188, 
    -314.785392363955, 
    -312.770576353169, 
    -319.474379997638, 
    -351.590921177709, 
    -409.212447551971, 
    -497.586514856353, 
    -562.663188699379, 
    -534.686652141881, 
    -297.691112441414, 
    -159.78764596151, 
    -107.614100715748, 
    -117.80947517254, 
    -54.3092457311012, 
    -17.7541756137355,
  
    -582.572252493556, 
    -228.639514957271, 
    -168.172831570581, 
    -141.72679506838, 
    -101.071870845483, 
    -66.5828322066706, 
    -47.8345205087011, 
    243.129118418508, 
    649.772743122575, 
    756.355956706598, 
    1532.69087058619, 
    1133.58783199059, 
    687.846018245482, 
    1022.69135464693, 
    906.854175571899, 
    797.228037177382, 
    593.743489196026, 
    614.136583753289, 
    651.845206018258, 
    527.187318607514, 
    382.098474867801, 
    281.87268755444, 
    265.801053300284, 
    228.396534914399, 
    232.383276726871, 
    231.678851248302, 
    154.134263389989, 
    145.659487624986, 
    139.220270075696, 
    138.592376358698, 
    143.953593297875, 
    328.564764323988, 
    382.910649554859, 
    201.320956214144, 
    233.522376458829, 
    221.454288217815, 
    214.61147832283, 
    118.171213290993, 
    223.9938137016, 
    360.293517694762, 
    524.49477848681, 
    805.790169522584, 
    1095.67849292307, 
    1440.58150271152, 
    1371.62899947728, 
    2573.54734687763, 
    2491.67763817457, 
    2096.18238668239, 
    1786.73729130829, 
    1756.70504039666, 
    1306.74412818558, 
    569.639668514847, 
    -114.139274062129, 
    -259.656821832946, 
    -352.844738925024, 
    -392.618447208725, 
    -336.620691827002, 
    -360.489664695031, 
    -493.870677251698, 
    -454.81599242583, 
    -353.943650723037, 
    -301.027331622424, 
    -315.201756134546, 
    -316.91736544687, 
    -327.994270123934, 
    -349.287982598932, 
    -381.984237995554, 
    -468.978047301495, 
    -519.183433443008, 
    -628.911027820754, 
    -440.658031805362, 
    -168.123810397551, 
    -115.061438099134, 
    -84.1571582802732, 
    -66.6223549832149, 
    -31.0382140056551,
  
    -528.499989350458, 
    -194.070758183085, 
    -206.538029697414, 
    -195.940275384491, 
    -134.24160708185, 
    -55.512867374356, 
    -48.3478595166564, 
    265.160541662579, 
    862.701344694031, 
    1174.49090673568, 
    439.469097598804, 
    700.730117182717, 
    635.509220785417, 
    564.647439407741, 
    577.977237492099, 
    504.028568378889, 
    523.948615139303, 
    517.991312682695, 
    363.398061609215, 
    359.790141892727, 
    303.241086150337, 
    292.912099695152, 
    217.173353150337, 
    221.578036544304, 
    221.978360439869, 
    168.486044175681, 
    133.784273865242, 
    131.588889898405, 
    176.546124843841, 
    124.271981248931, 
    185.630764050286, 
    172.91221430267, 
    265.919891457808, 
    184.194056441509, 
    181.892524413807, 
    202.891785060972, 
    98.8527086616766, 
    129.717795840839, 
    363.659275426577, 
    336.488993906362, 
    594.452812733068, 
    857.387633431534, 
    1258.96985562144, 
    1718.96181640967, 
    1695.4611236128, 
    2080.76587377124, 
    2385.04910476531, 
    2229.55294280357, 
    2554.83875266969, 
    2185.00955340309, 
    1665.96117658284, 
    940.21189422436, 
    46.3082010374849, 
    -215.060221754291, 
    -395.215155841789, 
    -365.563583121988, 
    -269.920278769191, 
    -299.790586375443, 
    -500.147293278779, 
    -455.915770958945, 
    -320.320050144515, 
    -303.050005986469, 
    -306.806413251102, 
    -309.634916166709, 
    -312.940545217721, 
    -336.927552841545, 
    -398.831914455333, 
    -475.95396543804, 
    -539.086869106314, 
    -661.025062279099, 
    -675.714278747625, 
    -340.28883928254, 
    -138.571134103773, 
    -100.002435642554, 
    -105.537559405687, 
    -105.242094253506,
  
    -533.371812608981, 
    -159.574479853853, 
    -186.612599391019, 
    -200.187345404374, 
    -234.249583753733, 
    -338.968515799801, 
    -202.394555453891, 
    -39.0751190282994, 
    240.770815203197, 
    618.875727065068, 
    415.988818596887, 
    403.445897622444, 
    166.642335023485, 
    373.29566930363, 
    330.2782872404, 
    260.362716873443, 
    402.989928639616, 
    320.747851603509, 
    289.619974779255, 
    306.77803684162, 
    233.41912087401, 
    261.673668217419, 
    275.691806370307, 
    205.333696933503, 
    186.992065835506, 
    136.789240924668, 
    116.18061066635, 
    135.130408881893, 
    165.931246331398, 
    120.840576590509, 
    184.308625863087, 
    119.026727423289, 
    261.022507927052, 
    190.167466267226, 
    121.371590117725, 
    109.799767887205, 
    99.6277797363639, 
    155.978669391902, 
    267.365638470196, 
    420.933640333735, 
    346.60733530316, 
    653.705333218464, 
    1165.11341493101, 
    1783.1529333749, 
    1974.20725544997, 
    2111.12165357498, 
    2350.40833008223, 
    2084.77654704642, 
    2237.63790121217, 
    2222.07062898745, 
    1761.16698255037, 
    1015.54270033713, 
    307.88999953702, 
    -157.324903904658, 
    -270.479454783817, 
    -211.640490569299, 
    -234.791557600358, 
    -369.151257398548, 
    -597.833779363857, 
    -424.119835796974, 
    -239.67879101624, 
    -272.765824722683, 
    -290.57269406292, 
    -318.954713234042, 
    -337.380124185013, 
    -355.193620196916, 
    -402.125314509615, 
    -514.183264195185, 
    -596.573543040243, 
    -674.977235672322, 
    -818.276948653304, 
    -595.169373635081, 
    -174.647291711035, 
    -112.211336028002, 
    -151.003301834073, 
    -114.091156654102,
  
    -582.842344166584, 
    -219.097189246474, 
    -170.185890212705, 
    -165.656658736482, 
    -118.857790736575, 
    -63.2894343347326, 
    -255.086980800479, 
    -265.242645084257, 
    48.9074464858841, 
    141.709222022523, 
    203.640402246029, 
    378.940914350555, 
    330.535375148692, 
    292.879693777804, 
    267.092205884876, 
    272.441487823862, 
    222.318342247308, 
    181.219464115172, 
    219.006135056294, 
    301.832588191529, 
    245.143195317814, 
    277.80863816367, 
    298.024598449502, 
    249.046417827969, 
    184.893728886313, 
    139.494865220979, 
    121.304258588981, 
    161.535463785938, 
    165.596337338711, 
    174.493354207858, 
    181.53027991565, 
    143.988072310957, 
    153.085286927517, 
    124.825100440594, 
    59.255013379378, 
    181.289459728313, 
    220.264558437557, 
    287.004604929105, 
    232.432270470819, 
    175.085354842371, 
    221.345214339681, 
    234.20135724024, 
    742.630804841492, 
    1308.13398189054, 
    1673.29432849094, 
    1821.35988826261, 
    1913.02983019787, 
    1945.44252079091, 
    2076.76351019677, 
    2088.21820488702, 
    1697.06563734714, 
    1097.763352534, 
    288.673512396855, 
    -118.627364017662, 
    -176.853329693751, 
    -196.788460657818, 
    -304.447935725915, 
    -543.991083356595, 
    -599.271836429267, 
    -272.582078929443, 
    -196.518532200864, 
    -256.017259497392, 
    -288.689732144688, 
    -310.719014897192, 
    -321.178078710165, 
    -339.88683545496, 
    -372.165001970656, 
    -511.230779487636, 
    -584.844758677724, 
    -740.811843444893, 
    -931.143085005572, 
    -776.719166216364, 
    -247.130926800734, 
    -177.173894971909, 
    -124.883874480962, 
    -88.9919150535097,
  
    -624.408482524876, 
    -366.987871236258, 
    -166.712245610099, 
    -131.168640925929, 
    -85.9866418913257, 
    -51.3493098838865, 
    -40.7723512136922, 
    -135.37653310355, 
    246.235119624206, 
    340.246402578151, 
    546.959067807085, 
    676.586976652584, 
    635.198431751896, 
    367.069348065077, 
    447.526274088383, 
    338.216299012153, 
    387.840695896981, 
    415.530878180219, 
    294.391398926465, 
    296.0615309601, 
    308.035375772371, 
    298.97325847237, 
    291.2074160688, 
    232.423195081755, 
    178.68932658, 
    104.702145152503, 
    79.9965921687119, 
    161.941962537947, 
    167.663018733897, 
    181.108230862078, 
    180.94142467204, 
    134.484277430467, 
    116.567838241646, 
    199.12409694411, 
    78.1842496856997, 
    191.467031286652, 
    279.300807256582, 
    411.380013191419, 
    157.110298733428, 
    53.1081397338515, 
    108.933450297305, 
    67.5457041485182, 
    532.289031952522, 
    924.216615239023, 
    1337.54425260709, 
    1481.46071485496, 
    1635.19278842631, 
    1727.39802875925, 
    1416.13124615882, 
    1593.50196701682, 
    1622.01721353734, 
    1198.55414139597, 
    477.295594820913, 
    -38.1033074839789, 
    -125.620655461362, 
    -187.478446135997, 
    -352.496764286637, 
    -501.376409562678, 
    -468.191914437732, 
    -185.984042544648, 
    -178.254773721984, 
    -205.627601926832, 
    -247.621688810735, 
    -285.125604084865, 
    -302.515115415396, 
    -324.865218492532, 
    -346.864379476994, 
    -500.627958086278, 
    -666.104654318542, 
    -830.657370905862, 
    -1068.25442829538, 
    -942.125988369693, 
    -482.522126952851, 
    -228.895411103729, 
    -177.407798572724, 
    -171.629991373316,
  
    -652.940084322836, 
    -497.743979237249, 
    -166.578824800446, 
    -107.084251099444, 
    -93.8728386023544, 
    -55.5895603474683, 
    -80.4424647622786, 
    -51.5329209518058, 
    443.522910435282, 
    622.238523929677, 
    972.487515550978, 
    991.006324657, 
    764.767890938718, 
    282.244076988333, 
    507.146714102647, 
    422.584157185485, 
    500.538200771421, 
    589.665635317197, 
    455.931637446797, 
    352.231668175401, 
    313.387315568572, 
    313.857869693974, 
    261.305407785755, 
    178.727599796496, 
    45.491247249744, 
    99.1555168092051, 
    -29.7529387949296, 
    163.051632499909, 
    112.428780758634, 
    69.7975400815749, 
    94.6953600630384, 
    146.191529621069, 
    177.997754783673, 
    57.2165673015366, 
    -22.7387917013743, 
    96.1749454019855, 
    187.671469614727, 
    231.9021342065, 
    152.826696348884, 
    115.149480687277, 
    127.090405168352, 
    239.586658804575, 
    486.904209085703, 
    406.792717112405, 
    1015.85144813598, 
    1401.92778684951, 
    2026.87846581266, 
    2009.52206161174, 
    1555.12198410803, 
    1455.83697819042, 
    1728.20918777996, 
    1386.51543692218, 
    912.218373177963, 
    487.933099381467, 
    -58.6082092885347, 
    -215.288185809523, 
    -434.980044459978, 
    -462.33900797247, 
    -406.928940686506, 
    -274.486171882603, 
    -215.222072464621, 
    -202.927127699302, 
    -246.620438102646, 
    -294.61814514707, 
    -295.941982192395, 
    -312.554609172689, 
    -303.776213625644, 
    -384.828526102816, 
    -725.476334455433, 
    -938.815261857909, 
    -1216.69618751381, 
    -1109.67436530956, 
    -808.373428532684, 
    -365.804816533308, 
    -228.098730928821, 
    -246.844692354106,
  
    -729.09469289235, 
    -554.590088257999, 
    -179.889413662747, 
    -101.944427999644, 
    -100.610358967626, 
    -56.8846073823439, 
    -53.3985349178848, 
    -55.0403209869965, 
    149.451100226611, 
    525.894245391198, 
    627.570783574529, 
    379.336852612983, 
    359.571095713309, 
    494.552726023676, 
    434.477117241563, 
    312.194235337143, 
    512.913138830649, 
    549.470641175684, 
    491.455299001525, 
    276.66878440105, 
    170.127838753104, 
    204.534997055805, 
    188.669884159477, 
    174.508919872869, 
    174.256256727195, 
    106.821894119194, 
    38.9923088617316, 
    70.685057520466, 
    64.7306374083173, 
    -22.6918744000984, 
    63.6564756854784, 
    157.995954686557, 
    122.252912643108, 
    137.573216659358, 
    -11.4425742991962, 
    41.2606136681384, 
    24.6604606662723, 
    43.6463829581971, 
    39.9895001867778, 
    212.80524442017, 
    178.377978575858, 
    440.399154440954, 
    373.234633387005, 
    504.40899833346, 
    863.84208146936, 
    1290.62458148542, 
    1731.31518522222, 
    2003.91310314422, 
    2030.94746855152, 
    2071.592514021, 
    1804.96210993204, 
    1740.9820121432, 
    1478.92788228102, 
    966.950003646388, 
    132.634798643703, 
    -148.687028209951, 
    -467.120583964621, 
    -379.05571753661, 
    -283.80917946195, 
    -293.0317278752, 
    -275.064796353775, 
    -246.104331799344, 
    -293.077527720076, 
    -266.327490269403, 
    -275.282206438156, 
    -269.905561496269, 
    -298.684153374205, 
    -309.004838599603, 
    -678.086243316548, 
    -896.666299134328, 
    -1330.57224281371, 
    -1174.36150830857, 
    -878.322440374871, 
    -512.688881962723, 
    -313.64759376842, 
    -252.10670225137,
  
    -774.647098220876, 
    -454.041797031347, 
    -182.09633543777, 
    -105.681717199815, 
    -87.4929653703833, 
    -50.7172263525635, 
    -49.9056345586147, 
    -47.3061528729164, 
    -41.4872168239805, 
    245.469542401901, 
    355.14496805633, 
    240.903632899814, 
    502.045866108688, 
    161.280901181602, 
    128.414762785293, 
    353.705458116691, 
    290.889412370535, 
    449.258837713774, 
    476.665691546603, 
    269.325041780546, 
    149.820518010941, 
    172.950264380733, 
    93.3409616602766, 
    173.496291200097, 
    104.086209290772, 
    95.2921638584883, 
    63.5103182632472, 
    51.6705305525597, 
    52.0346044276623, 
    11.7857190647558, 
    22.263738730186, 
    46.9174940481961, 
    30.9009415657496, 
    100.464486260964, 
    -13.502564885582, 
    58.1602619108137, 
    50.3284019606912, 
    20.64267487889, 
    -88.1159892514735, 
    174.597230966789, 
    308.889184659166, 
    384.431638288338, 
    382.52493957229, 
    530.547342904871, 
    752.779416330986, 
    993.76402326287, 
    1184.34405086983, 
    1597.56177699312, 
    1754.16459454134, 
    2007.45395818456, 
    1905.96439628986, 
    1696.87511185223, 
    1724.62376909587, 
    1129.85728251253, 
    689.968774015932, 
    -250.794742413366, 
    -234.961658655059, 
    -165.00123019715, 
    -187.509889414703, 
    -247.027916954186, 
    -301.014577457646, 
    -295.361006780541, 
    -264.719742756808, 
    -267.983441274884, 
    -241.720701657644, 
    -280.175018082008, 
    -337.699541700647, 
    -318.721221611988, 
    -442.957589233844, 
    -976.039528063941, 
    -1385.21564137629, 
    -1250.18462367554, 
    -970.594586994987, 
    -684.18564036712, 
    -471.730365155124, 
    -360.53125641621,
  
    -648.790348928691, 
    -263.759994079658, 
    -179.609547537091, 
    -120.851886705482, 
    -98.8461282853985, 
    -51.7301741020143, 
    -46.943176370986, 
    -33.0392327858646, 
    -55.6473484461146, 
    130.205952725511, 
    151.634558493988, 
    132.357995959171, 
    228.578666330319, 
    238.946924034452, 
    146.141529886344, 
    177.985999866669, 
    186.784058759888, 
    452.923962545021, 
    369.011039281077, 
    290.931658792869, 
    67.4201630526111, 
    -6.13222457486863, 
    112.559846284275, 
    77.67092486218, 
    5.1391258554773, 
    46.4203153412125, 
    76.7213562851123, 
    56.9413601169392, 
    42.7558499397116, 
    31.5077575660098, 
    -45.3086652857198, 
    -51.7589462073097, 
    -12.2674146250541, 
    69.5619026442523, 
    44.3343190356573, 
    1.15996145921681, 
    -43.2788524566275, 
    -35.3217965384485, 
    -74.7051734262191, 
    128.76205882567, 
    332.217046103312, 
    364.606530701058, 
    256.270494206887, 
    469.129205859656, 
    618.700307156177, 
    941.160290973318, 
    1259.28207441887, 
    1338.31438072692, 
    1669.68564102498, 
    1918.46935903586, 
    1914.78881157579, 
    1257.95711615586, 
    1683.30452143038, 
    1084.32842766397, 
    340.520633398488, 
    269.857440884425, 
    368.12154791684, 
    434.163492422761, 
    188.063368569833, 
    -63.247017188473, 
    -333.584387126722, 
    -294.039973242952, 
    -277.75791620167, 
    -333.682307411016, 
    -357.976084556453, 
    -392.541690151476, 
    -322.033920125758, 
    -313.886543329459, 
    -457.772305713924, 
    -1090.40990283962, 
    -1367.19524888469, 
    -1408.53744783647, 
    -1109.22767849332, 
    -846.672714549509, 
    -532.315027008394, 
    -514.951655986996,
  
    -324.472628765382, 
    -212.946651181075, 
    -192.049826230074, 
    -143.38239443182, 
    -106.741685303435, 
    -54.9156099497805, 
    -37.0755057110631, 
    -30.0723051699119, 
    -91.0503169302179, 
    33.5746821291897, 
    124.867178351988, 
    213.630889572194, 
    141.748100022319, 
    214.79699613052, 
    199.61126234176, 
    169.17974413309, 
    289.749432188933, 
    413.651889848015, 
    391.200652320068, 
    103.065243707657, 
    34.0332394233613, 
    99.941333001833, 
    62.8429129646987, 
    67.5659876804206, 
    13.2749642259873, 
    58.2489643277125, 
    87.431030101499, 
    29.2028108656916, 
    0.895168294297731, 
    57.7005081784055, 
    -153.973486837321, 
    -140.614467462794, 
    -103.153584576401, 
    37.0130835270958, 
    185.894639206359, 
    -60.2626815744647, 
    -95.9343089074861, 
    -72.2415284843486, 
    -48.711871862678, 
    76.8448326320698, 
    144.033424665784, 
    177.020490917619, 
    219.449594200793, 
    369.747024228565, 
    416.256842033326, 
    585.107144841689, 
    495.918344674953, 
    1103.67082344217, 
    1173.73658185149, 
    1454.28463203455, 
    1726.92238059049, 
    1493.54312824108, 
    1468.36002531831, 
    1217.34626182223, 
    233.758346047144, 
    1120.04091865566, 
    951.735940042566, 
    518.500066152749, 
    498.724378562322, 
    89.3339210388868, 
    195.396458250143, 
    -159.124032709392, 
    -221.723655929223, 
    -500.893826808267, 
    -413.557868457718, 
    -261.744553218895, 
    -243.084140858751, 
    -327.173817317404, 
    -492.982415757815, 
    -1140.90192347545, 
    -1421.17219787803, 
    -1472.27509045574, 
    -1298.93678681821, 
    -1013.2967146631, 
    -747.283718677277, 
    -657.197493515784,
  
    -232.923471457213, 
    -212.543928063063, 
    -202.255807778336, 
    -159.805498445688, 
    -115.473237262995, 
    -79.4959461750401, 
    -42.3957796812327, 
    -32.15473682536, 
    -123.668025741919, 
    -19.4664372408664, 
    73.8687481186023, 
    155.533938045864, 
    90.8788865037073, 
    133.036946768723, 
    29.283566351301, 
    278.096519809819, 
    248.227175824721, 
    302.328559772965, 
    216.044897697804, 
    110.072263843134, 
    131.998697244576, 
    205.48886943531, 
    175.67121442515, 
    8.42633088508703, 
    -44.5374252688077, 
    -334.145033307734, 
    -20.9650968206788, 
    -86.6528960678635, 
    -53.5042797555307, 
    -47.5551204029953, 
    -48.7336717757232, 
    -143.49678223344, 
    -171.559690080324, 
    -139.618869869066, 
    -78.5262283461903, 
    -60.106046475994, 
    8.25238338997321, 
    7.29436404866298, 
    26.0693896027727, 
    68.701498805342, 
    125.018633296749, 
    170.442174986256, 
    310.720274400872, 
    391.56488442501, 
    363.915434898215, 
    228.014335194465, 
    234.723985603651, 
    853.40560474802, 
    914.376442023916, 
    1443.69249837262, 
    1644.60455259043, 
    1216.02636663216, 
    1060.56325115787, 
    430.705471478826, 
    1409.42283650875, 
    1617.08722038311, 
    1597.91446353447, 
    1081.07834075894, 
    32.0211086764277, 
    280.339838134767, 
    699.265764546144, 
    322.37410220267, 
    -72.923209441335, 
    -219.750575167066, 
    -227.2397970112, 
    -186.366224835728, 
    -256.252988612399, 
    -299.836799583136, 
    -414.816747005417, 
    -943.165278871546, 
    -1358.83943183104, 
    -1459.4406964002, 
    -1435.95192832135, 
    -1203.1345238424, 
    -968.391786410854, 
    -775.450625976017,
  
    -277.342241712274, 
    -270.439428686162, 
    -237.166488504357, 
    -168.547659172323, 
    -138.690534862933, 
    -97.4190923620312, 
    -55.1168972855854, 
    -43.8977215821375, 
    -249.140003693464, 
    -145.051242829638, 
    10.6713086990065, 
    72.3857090182162, 
    147.193662940323, 
    194.158363098795, 
    104.201589874834, 
    154.855012266795, 
    324.929653496651, 
    310.28740029586, 
    -21.1571274638699, 
    -74.8280160269566, 
    104.900244640208, 
    140.620449461302, 
    116.892916187058, 
    76.2703308092658, 
    36.6163241084893, 
    -108.291528027907, 
    -153.073739711806, 
    13.7781685004724, 
    6.14581119760473, 
    -46.0772365127414, 
    -145.251202946414, 
    -48.4574076432522, 
    -61.1903959885147, 
    -89.8775517345139, 
    32.1390854311173, 
    120.747777519141, 
    120.274765620173, 
    37.1829488878151, 
    115.340622221637, 
    39.1489054620058, 
    97.8785206665517, 
    227.847859584471, 
    314.816848985559, 
    363.684620813453, 
    339.727561356905, 
    195.179355044651, 
    448.101598199246, 
    1048.06047480157, 
    1369.36140694784, 
    1339.11132595494, 
    961.400343917382, 
    666.534539986294, 
    398.774081517441, 
    1180.33667298902, 
    1934.75661551379, 
    1848.35963164839, 
    1770.801599415, 
    739.900515271185, 
    705.774380366741, 
    1117.46159921543, 
    1070.92413141265, 
    1293.62749957077, 
    390.228753541653, 
    145.388667894246, 
    -129.119071456378, 
    -244.962882418918, 
    -294.655820237828, 
    -304.052949420549, 
    -309.262601863097, 
    -831.606337697886, 
    -1251.40426239321, 
    -1445.20673738588, 
    -1439.30398163149, 
    -1302.73398900219, 
    -1120.78182270866, 
    -912.726956503123,
  
    -320.99193587095, 
    -316.819878209746, 
    -280.41149667396, 
    -197.218538895166, 
    -172.389780634062, 
    -157.37458695116, 
    -205.010903951173, 
    -280.228491105002, 
    -249.932647482946, 
    -375.152835115476, 
    -26.7256924566765, 
    84.8418074257562, 
    72.2901374116332, 
    219.688793404503, 
    -18.9978369949675, 
    43.8309901251893, 
    278.473839453328, 
    275.383358390439, 
    118.078256707445, 
    202.044267355397, 
    -20.1700852979876, 
    128.005144387048, 
    -128.984811524396, 
    116.638897495334, 
    131.982556801227, 
    139.588096963597, 
    54.2402714198545, 
    209.603843385667, 
    13.3774600561636, 
    -61.0821498639104, 
    -90.6051654997215, 
    -18.075392606678, 
    -100.397074815811, 
    -172.396880932645, 
    -26.475154696227, 
    -31.9960046909186, 
    1.09810511796105, 
    69.5401148673274, 
    96.7924505791219, 
    -23.80171649213, 
    121.728069035232, 
    226.116676821822, 
    279.170557831597, 
    377.122113064449, 
    421.985753472683, 
    536.177948245814, 
    842.473242397676, 
    1140.6276745086, 
    1438.11811406561, 
    1255.14132977492, 
    991.052887313177, 
    929.15768823912, 
    730.737585420179, 
    1943.8970183301, 
    2183.09745431454, 
    2109.35220374506, 
    2183.51674519675, 
    884.732624852785, 
    1568.15941882161, 
    1865.87836971478, 
    2293.66559900708, 
    1308.73580141483, 
    1160.12468038561, 
    876.552820254815, 
    406.448481313068, 
    -106.78007467303, 
    -245.409443794412, 
    -286.677880290373, 
    -249.862019031606, 
    -369.473251171901, 
    -1007.43599570212, 
    -1395.44614756414, 
    -1478.630559257, 
    -1400.12916582029, 
    -1266.20691251167, 
    -1032.33905364204,
  
    -398.708587172317, 
    -379.205874704701, 
    -374.806830898512, 
    -326.874365551343, 
    -358.87264061188, 
    -480.772347829378, 
    -485.740644123892, 
    -426.778744064279, 
    -290.645549120588, 
    -613.205943980114, 
    -215.017076060863, 
    -24.1131352682846, 
    66.1634236140321, 
    3.24758602002847, 
    -200.105904328196, 
    -10.4987923930795, 
    199.514987189455, 
    149.279566257558, 
    339.629059331283, 
    252.783803997488, 
    62.4316286944592, 
    83.8569092168477, 
    122.219130180715, 
    22.7206579461457, 
    112.803858783716, 
    21.0845923031615, 
    -15.4020399760221, 
    -11.89733014809, 
    33.8607709559986, 
    -11.87500380315, 
    -76.4023391023066, 
    -41.8274009657602, 
    -86.6138019326822, 
    -147.451027644841, 
    -113.472097181126, 
    -184.162277640312, 
    -105.095672513174, 
    110.181836336483, 
    -3.92880628764528, 
    24.6364729834301, 
    35.4951743035675, 
    126.160280024751, 
    243.961851141355, 
    436.758905246303, 
    523.659985626666, 
    724.840062644422, 
    1037.75684538667, 
    892.227017179447, 
    767.449099627211, 
    656.478584562947, 
    1103.16548178952, 
    894.485614396427, 
    1386.84701777307, 
    2161.95494908315, 
    2384.74936446204, 
    2296.62838789544, 
    2380.76371493452, 
    1732.30546650134, 
    1599.46071511127, 
    2122.23880384216, 
    1916.08658604125, 
    1591.64989151053, 
    2164.86979068699, 
    1588.94345603678, 
    990.292453624901, 
    755.623897274827, 
    78.4795719562713, 
    -146.734210688215, 
    -279.310087308637, 
    -315.431609244524, 
    -719.004942907862, 
    -1145.47438977146, 
    -1434.65341160893, 
    -1483.76464602822, 
    -1312.33964309607, 
    -1139.44077042156,
  
    -328.740722118005, 
    -342.658027290095, 
    -339.161139331232, 
    -364.908144050589, 
    -391.233031218422, 
    -448.010564831842, 
    -349.767006834569, 
    -352.354554798939, 
    -297.072860798937, 
    -355.379604988904, 
    -795.36398506805, 
    -330.589557472569, 
    -364.920050143661, 
    -237.515467849853, 
    -130.051022182523, 
    -268.45539219035, 
    205.438268473539, 
    98.4446757477858, 
    267.1593537966, 
    -186.70921738553, 
    -115.13872149814, 
    47.3308955883389, 
    -168.887203501703, 
    32.2109001132742, 
    129.096296761099, 
    -89.3034995934466, 
    -69.8934596863732, 
    -94.381364299095, 
    -23.6420879484517, 
    -71.8097933815161, 
    -176.347349549194, 
    -134.432357983521, 
    -43.8749216724199, 
    -63.6158236453405, 
    -66.2768845782427, 
    -50.0060942944584, 
    -42.1935600855303, 
    53.9177667333729, 
    51.4563806903333, 
    28.9999724101904, 
    51.7176014210327, 
    204.349047497433, 
    260.425050985373, 
    389.717366255945, 
    470.268537019428, 
    681.084498748267, 
    948.737186675376, 
    781.653551142268, 
    885.699460088344, 
    1203.6614505644, 
    1347.09812469311, 
    1050.51919956356, 
    1366.98900174507, 
    1754.6651554428, 
    2260.08877085037, 
    2542.58352350148, 
    2382.66770605277, 
    1966.90710478267, 
    1626.10415919391, 
    2240.7827051041, 
    2064.38952689688, 
    1877.49429056439, 
    1631.29735572875, 
    2050.79032715117, 
    910.304061667521, 
    1255.41854569627, 
    628.130623513083, 
    -9.04594356121974, 
    -260.147636607941, 
    -231.833081979099, 
    -250.876957420273, 
    -312.432418801883, 
    -1324.31181441389, 
    -1452.34356450234, 
    -1412.20813439381, 
    -1236.72778783373,
  
    -330.21515051061, 
    -324.485313257472, 
    -349.95186328354, 
    -352.960889762887, 
    -343.036538904752, 
    -325.609650990998, 
    -201.450475876438, 
    -247.137149052551, 
    -229.478180266973, 
    -170.23124755697, 
    -211.94096120982, 
    -395.962635625529, 
    -290.137040927451, 
    -352.893860640741, 
    -371.448293623969, 
    -310.587904961085, 
    -165.121004623902, 
    -252.040377279427, 
    8.62474827582339, 
    -33.1638194342613, 
    18.6523077338387, 
    124.882583790098, 
    -50.9039899985246, 
    38.6542564989267, 
    -10.5129931299756, 
    70.6419349984886, 
    13.1786567865117, 
    -218.746046012884, 
    -193.032967993554, 
    -129.141150960465, 
    -124.595528344158, 
    -80.149737444598, 
    -9.34617089939877, 
    -4.61718062377407, 
    -22.0629808177221, 
    29.3135808344503, 
    45.4279527904464, 
    -35.3917732842124, 
    23.7345220121561, 
    -14.496258677854, 
    113.774855986421, 
    170.688461709531, 
    199.020510347802, 
    281.118402013322, 
    262.297829340716, 
    523.325780712614, 
    819.005711955964, 
    949.935450939425, 
    1283.53581261715, 
    1333.49431898025, 
    1250.51508513276, 
    1089.76648289252, 
    1181.94626766944, 
    1495.10467787313, 
    1844.45413491655, 
    2099.09909153306, 
    2271.46872723997, 
    1939.44215261495, 
    2023.24459673121, 
    2055.87411068428, 
    2152.16684472574, 
    2377.88748473095, 
    2408.1111711628, 
    2595.43743028459, 
    1916.41917231474, 
    1764.50473099353, 
    1197.25792970048, 
    235.154045151958, 
    -114.480724083219, 
    -317.635802111991, 
    -357.258978246707, 
    -308.662504856157, 
    -1029.11603668316, 
    -1492.41966931043, 
    -1472.65268427901, 
    -1464.54763269371,
  
    -331.589859781981, 
    -320.609765726668, 
    -306.47384211678, 
    -315.54179982509, 
    -289.662114266186, 
    -186.224441872198, 
    -137.662901676515, 
    -162.338758767653, 
    -200.94168761703, 
    -151.086093293859, 
    -105.018181780552, 
    -295.319240834917, 
    -553.571507350329, 
    -490.610703480071, 
    -368.110055652205, 
    -306.538510295873, 
    -269.79751458333, 
    399.845020618843, 
    -9.61496075377262, 
    135.12446076712, 
    262.379759337845, 
    248.018665918178, 
    221.527126243906, 
    150.708749762576, 
    -33.2907936682464, 
    49.2428974875699, 
    77.922753875492, 
    -126.636952725934, 
    46.7517802766021, 
    34.1212733289822, 
    26.4139247549329, 
    -47.2079396811195, 
    20.0134632488646, 
    47.5311282297795, 
    65.4271999585533, 
    136.166946525404, 
    56.7482926284883, 
    -145.304899249874, 
    -136.877535241182, 
    -72.2235259203468, 
    64.393908667673, 
    73.3498417858587, 
    76.6626308655833, 
    104.490651099707, 
    149.877798286559, 
    320.536527302607, 
    573.912122634602, 
    732.361420976359, 
    1410.66116572227, 
    1193.42719402933, 
    1094.53636036155, 
    1031.39143720159, 
    1002.37967139369, 
    1281.29731875225, 
    1410.47546383301, 
    1839.65551715095, 
    2266.52429558049, 
    2338.25767320588, 
    2361.93626682328, 
    2473.20392970035, 
    2395.96091583355, 
    2478.68216755729, 
    2309.60576052949, 
    2369.96956238956, 
    2101.31096610724, 
    1777.9089141709, 
    1202.5750709696, 
    451.311410918884, 
    44.1656315113756, 
    -266.225658734998, 
    -220.713116230384, 
    -305.537801740418, 
    -1042.88945372134, 
    -1263.87012164724, 
    -1343.8814589446, 
    -1392.22937382509,
  
    -343.141554367902, 
    -316.902398774765, 
    -300.050006054817, 
    -297.402986310765, 
    -244.154100031495, 
    -198.099269751605, 
    -151.40260274573, 
    -151.763330119989, 
    -168.583573598745, 
    -133.442785709462, 
    -150.30946782562, 
    527.839045670902, 
    303.598693418332, 
    49.9486900812149, 
    -198.415320135952, 
    -264.099625026794, 
    -141.925955769203, 
    246.154827986156, 
    402.134098206758, 
    364.858872066552, 
    160.856011054277, 
    215.120197157311, 
    283.439994397647, 
    136.127819836608, 
    -13.6816141329313, 
    13.0817286354492, 
    14.3413551724782, 
    33.879857949153, 
    74.1390349611331, 
    -81.3297289830183, 
    -73.5439012501836, 
    -33.989178125228, 
    30.045420413055, 
    77.1918937772813, 
    62.8323439686725, 
    16.9135148300993, 
    36.3155636557146, 
    -34.8421067235719, 
    -47.6859809196282, 
    32.552694524389, 
    36.9116252533935, 
    24.0567244783895, 
    17.9546115494519, 
    -9.31043732193123, 
    13.3376192814977, 
    215.007928929432, 
    335.770903084341, 
    628.64008152739, 
    961.967518634524, 
    946.0088770184, 
    794.773465779168, 
    800.597949746743, 
    931.543367810908, 
    1226.48965592507, 
    1393.3692063762, 
    1701.99599368789, 
    1967.22713221843, 
    2317.79985659814, 
    2427.94979345785, 
    2415.74001955585, 
    2426.70539686794, 
    2241.61141448325, 
    2082.6799405601, 
    1957.70262721832, 
    1887.74588016113, 
    1702.06116648777, 
    1331.3814021983, 
    836.942882226004, 
    651.990434952039, 
    -115.644585835849, 
    -184.501576441801, 
    -266.804232534343, 
    -502.965881616785, 
    -625.836840271824, 
    -589.148668252885, 
    -847.355145453348,
  
    -424.525059446907, 
    -320.062897903255, 
    -303.334502234037, 
    -285.564025426098, 
    -238.919575335598, 
    -202.908342337955, 
    -163.794888149317, 
    -190.610287368364, 
    -213.31436641646, 
    -176.461716185226, 
    31.4328793902386, 
    147.828220745483, 
    407.006756089438, 
    965.671726179816, 
    564.833131420647, 
    -76.7853601115021, 
    83.444625794694, 
    123.922634058848, 
    192.029578338149, 
    165.252193405541, 
    209.683797031076, 
    376.327165498978, 
    391.09986614727, 
    216.031314941694, 
    153.306693460479, 
    112.660711256413, 
    -85.6567278196687, 
    -76.8552392581025, 
    33.0601574106417, 
    -59.1140785818018, 
    -84.7471427669194, 
    -12.6155736483848, 
    15.6786683078305, 
    87.8727879198495, 
    -25.1120773541832, 
    -80.9053887375804, 
    -23.9291827683683, 
    -86.6496825111396, 
    -19.5132200878115, 
    37.9276955872607, 
    32.699914260781, 
    18.7153322613921, 
    47.960156792089, 
    127.868777580519, 
    171.841660923545, 
    229.134302812087, 
    303.800682947858, 
    429.103534454996, 
    596.665757361881, 
    668.819878128583, 
    645.135272872941, 
    747.417728154951, 
    873.754912552617, 
    1224.01084802506, 
    1453.98934316261, 
    1203.163791413, 
    1448.73335043982, 
    1857.88342303953, 
    2234.25619728969, 
    1854.99884578283, 
    2163.19970979937, 
    1912.96936674214, 
    1913.84394641633, 
    1598.97954696878, 
    1652.42157672742, 
    1451.94941530303, 
    1199.72249457177, 
    1072.73402676471, 
    741.796405557283, 
    503.397155266183, 
    -199.205057789208, 
    -218.066596365455, 
    -253.814348161021, 
    -328.832886054028, 
    -362.914437972151, 
    -387.500213165967,
  
    -871.432040326666, 
    -440.887573947029, 
    -304.477212198905, 
    -296.730849754103, 
    -246.972259314303, 
    -200.103327884652, 
    -189.181968923912, 
    -242.036478181435, 
    -237.53674309358, 
    -107.683988429132, 
    415.5357076553, 
    502.739418196383, 
    789.738918090851, 
    1260.52644906893, 
    514.898072668843, 
    -249.237999359671, 
    -280.823906833354, 
    129.171033468396, 
    178.521407919798, 
    272.250800941184, 
    154.954292004745, 
    384.008110717057, 
    469.367220584917, 
    365.102233600509, 
    253.863300949301, 
    119.70566052739, 
    136.62390877872, 
    221.330632236476, 
    116.171248009864, 
    46.5072961670566, 
    96.7975795602742, 
    26.8676369361085, 
    53.8661621703548, 
    71.098595791141, 
    1.52244946260342, 
    0.699248184573447, 
    13.4969738875352, 
    -50.1076317484948, 
    -37.4999323168895, 
    8.85438311739965, 
    13.6388351196405, 
    -11.3571429639084, 
    39.0559196648385, 
    190.166423464409, 
    240.240229690996, 
    254.242912014814, 
    241.704424850617, 
    361.304560478697, 
    488.328471898232, 
    580.397165723505, 
    639.028578686688, 
    737.773018848723, 
    907.345336700476, 
    1087.77950296263, 
    1442.26818611854, 
    1624.2905335122, 
    1434.50831364784, 
    1665.26705510566, 
    1679.86353906032, 
    1619.57446974255, 
    1443.53971131465, 
    619.418085266998, 
    530.428820722185, 
    854.498694211615, 
    1537.73474678134, 
    1470.85745876606, 
    1772.71263479679, 
    1336.07522232721, 
    1045.48966580141, 
    835.801922250297, 
    140.577932751844, 
    -161.279486127558, 
    -233.745857211003, 
    -337.88541925394, 
    -395.768128953616, 
    -411.077580493615,
  
    -1374.81666296674, 
    -654.384337866292, 
    -353.823934450395, 
    -287.748270395755, 
    -245.973328033994, 
    -209.908441396203, 
    -221.094679043248, 
    -176.569316947314, 
    -112.112416687097, 
    8.78633206956217, 
    461.093777219762, 
    595.088100228307, 
    1059.9390227776, 
    1240.86666494201, 
    -362.831987169526, 
    -202.364901679099, 
    283.253386771954, 
    305.205041020334, 
    224.003218301599, 
    372.427351422966, 
    387.510423688046, 
    417.554362507443, 
    487.065222002225, 
    456.071105311994, 
    284.876627158478, 
    105.482394711835, 
    153.539655703581, 
    214.216653027168, 
    48.4452665765247, 
    -47.194954974653, 
    43.607203787948, 
    68.8266047673157, 
    49.0858518602064, 
    27.3219725435557, 
    61.9150584205937, 
    70.1670323822557, 
    72.5431418018401, 
    61.5932272134661, 
    -18.5407494079632, 
    -23.8447095277192, 
    -19.8776170911073, 
    -20.3048860452746, 
    8.87952208418902, 
    32.2257197223612, 
    227.860708646786, 
    244.523789434659, 
    343.862953258657, 
    406.111912341829, 
    472.857636933365, 
    538.941217164043, 
    627.385063701087, 
    704.423624053647, 
    830.657550482843, 
    1102.34434758749, 
    1374.68242131796, 
    1576.0842143675, 
    1401.12473639715, 
    1430.12598290182, 
    1046.18854850778, 
    1188.04146316205, 
    1184.02696648372, 
    280.515257071798, 
    -437.414974283142, 
    1339.95377773188, 
    1503.1352543847, 
    1637.25456895648, 
    1908.64932673028, 
    1745.74086699107, 
    1357.23934531558, 
    803.225517947882, 
    512.35921477416, 
    -57.8051799840139, 
    -246.786747967677, 
    -407.1144386881, 
    -419.260580000925, 
    -410.183601426385,
  
    -1420.6884805438, 
    -975.403925281623, 
    -391.209115202456, 
    -287.532192430998, 
    -249.684832191681, 
    -202.580134745274, 
    -191.353174038724, 
    -126.808456777592, 
    -98.8211471124032, 
    -95.1496237288128, 
    283.51155242835, 
    549.258059109703, 
    1093.76832842854, 
    1157.60580106012, 
    -367.051419808111, 
    359.403815018501, 
    851.518628068093, 
    812.89519375142, 
    576.320939212474, 
    505.845800278035, 
    364.647066989911, 
    384.495041004621, 
    517.806475802738, 
    367.655321712858, 
    272.788658881107, 
    192.475537463505, 
    181.491044603029, 
    162.428729333909, 
    -42.7376687222338, 
    -166.812077100439, 
    -67.0133220036101, 
    25.5396418785065, 
    4.97390967130212, 
    1.45254646842357, 
    -53.2901799537296, 
    -71.7418577177113, 
    73.99328923092, 
    99.8528068436743, 
    -70.3758683327465, 
    -50.1068657643315, 
    -31.8879995815964, 
    -3.03933417728672, 
    11.5861403521937, 
    53.9077823073974, 
    137.502788315162, 
    154.871563034656, 
    218.581225872574, 
    323.664291706492, 
    345.628590898846, 
    489.001437021664, 
    586.315680979081, 
    769.769564390449, 
    908.597547917725, 
    1061.62673138558, 
    1214.87941655654, 
    1439.74971457692, 
    1611.90087757345, 
    1354.78333385847, 
    1472.12872558799, 
    500.860961738937, 
    1509.09621281639, 
    1242.08090153576, 
    1272.93577522712, 
    165.169060861957, 
    80.4763939121747, 
    1405.75405919674, 
    1291.54540106591, 
    1379.90027057097, 
    1531.47698010896, 
    1212.92490891887, 
    967.456200312391, 
    67.2241450940621, 
    -331.777934190809, 
    -468.139677220737, 
    -415.611089131867, 
    -360.345397838153,
  
    -1315.1333435332, 
    -1044.47107793076, 
    -413.758622587061, 
    -311.970903206512, 
    -266.984392821855, 
    -213.67360200914, 
    -167.855712320343, 
    -151.583277818737, 
    -116.088428857212, 
    -84.5152450926762, 
    83.1453529296008, 
    1005.0350486781, 
    857.38672306023, 
    -348.130768580502, 
    577.688963158529, 
    502.766547618492, 
    1038.09897845056, 
    27.1777777794657, 
    119.493860791533, 
    376.681050295257, 
    466.455409226199, 
    350.328810872317, 
    382.241057238947, 
    363.221966639878, 
    315.923597842021, 
    202.88949630669, 
    189.012155891667, 
    175.816864084155, 
    -48.4313303511198, 
    -165.278043885782, 
    -31.7766946016211, 
    17.3979873825427, 
    20.328219958943, 
    37.108533581054, 
    -58.6601652196646, 
    -120.904671795023, 
    15.0186756196512, 
    -9.16032880497871, 
    -59.2921274816335, 
    -48.1536318238612, 
    -19.7176803164893, 
    10.6980837052238, 
    86.9786043428773, 
    87.224797308644, 
    126.733813184372, 
    162.713146814174, 
    165.407018533346, 
    312.060473421787, 
    389.983913763373, 
    401.19226130179, 
    517.24852909887, 
    775.937198062227, 
    872.694430531741, 
    954.697244129417, 
    1056.6157972842, 
    1272.54940720715, 
    1433.77428671227, 
    1449.10081264927, 
    1480.52895299692, 
    945.778814386272, 
    19.5419464714578, 
    596.39176957151, 
    69.3634019805635, 
    1133.84213503961, 
    -234.481781390867, 
    10.0264673713858, 
    223.437394304483, 
    576.121731974925, 
    70.2730864261115, 
    -233.690422805658, 
    -111.635346362454, 
    384.377275514988, 
    -83.2783196589243, 
    -481.297688248176, 
    -482.508644377397, 
    -349.708736176187,
  
    -1121.74765583649, 
    -698.613150234583, 
    -313.858885052756, 
    -305.741299098443, 
    -309.533203731593, 
    -279.002231081016, 
    -225.844538762349, 
    -151.920781580892, 
    -103.786853863972, 
    -86.8657152297647, 
    -212.674193039453, 
    -38.4240738874396, 
    -166.349250466655, 
    523.645676897993, 
    363.83878527617, 
    1376.22244604438, 
    -123.971087204805, 
    -135.337406086905, 
    102.377034364063, 
    486.389618428265, 
    527.173622981433, 
    303.819790377729, 
    429.051184398998, 
    391.192372308199, 
    311.967610845104, 
    133.441720915534, 
    119.115606653999, 
    246.321444802963, 
    164.272079224283, 
    22.7840152730609, 
    12.0407940515078, 
    29.7051421960557, 
    17.1160832863773, 
    -42.4769968335058, 
    -108.491091340546, 
    -74.6819429210679, 
    -72.2260951248287, 
    -65.0282935556865, 
    0.410455412355306, 
    34.7124326072918, 
    6.07202787905989, 
    87.5166735195238, 
    94.6675982192277, 
    167.346694568236, 
    244.570534318452, 
    174.352718735597, 
    212.673820692107, 
    348.702234308771, 
    378.372582959968, 
    419.405901145294, 
    509.274089945658, 
    528.070572326592, 
    688.154517144934, 
    802.595178021028, 
    972.758559403201, 
    1135.51277208489, 
    964.007602875337, 
    1744.67758012966, 
    1175.46464208792, 
    1583.53747353548, 
    1155.16407871565, 
    197.340659984176, 
    1440.53607498973, 
    1158.88627976506, 
    208.918631268514, 
    -563.132454388357, 
    -502.835500351929, 
    -529.754191220272, 
    -443.438808757272, 
    -393.507182976699, 
    -411.830376799135, 
    -514.004562758117, 
    -451.600448313648, 
    -551.150437640183, 
    -499.274044024047, 
    -331.375207275185,
  
    -699.906482282168, 
    -401.98143557712, 
    -309.903344725709, 
    -305.287483847555, 
    -344.369990627549, 
    -325.444121677959, 
    -281.027565570589, 
    -241.569165055723, 
    -146.483403815669, 
    -77.6972029259864, 
    -31.1732895638637, 
    -431.796084306808, 
    488.324722755665, 
    1349.87525495676, 
    1091.24306820382, 
    430.651088573082, 
    -309.326740585288, 
    -230.865847554486, 
    -122.781238267292, 
    515.877377000661, 
    606.812061758349, 
    410.295257260793, 
    442.719270490452, 
    275.973288131321, 
    229.36897256046, 
    23.2721319641809, 
    249.70383940779, 
    350.954999148378, 
    219.468064490785, 
    108.567829253826, 
    52.0541880341685, 
    7.31150552126552, 
    42.1431069027005, 
    -21.7711985760016, 
    -2.56818337493141, 
    16.0281027834475, 
    -8.31365903113949, 
    51.3590459236262, 
    162.824807371031, 
    133.204147413623, 
    106.107752239317, 
    124.21269518157, 
    118.452969161287, 
    147.564303332989, 
    255.444823157214, 
    218.122290230011, 
    281.087749434212, 
    352.350647216148, 
    262.662585503044, 
    384.357038201037, 
    589.157126423494, 
    579.173848125462, 
    635.022513813562, 
    730.775176532058, 
    979.995184878092, 
    1409.03258086373, 
    1332.86107750836, 
    1276.63345675239, 
    464.288722885169, 
    1180.3345355539, 
    756.809958843441, 
    702.471640713939, 
    984.060923466337, 
    1889.88608953427, 
    1172.24235367214, 
    296.186677234302, 
    -438.079363153335, 
    -325.026651034294, 
    -160.292909094088, 
    76.5268808858309, 
    123.350616920707, 
    -237.025299933024, 
    -353.804450470811, 
    -485.085241849584, 
    -373.750460031983, 
    -307.98548960926,
  
    -523.761562091105, 
    -471.333337969637, 
    -380.986209583177, 
    -321.321626554279, 
    -335.493186002349, 
    -376.382152429221, 
    -369.643734674572, 
    -307.044746608245, 
    -247.131379307989, 
    -166.827531895745, 
    -345.682134703054, 
    -268.90413561327, 
    711.393592125345, 
    329.377145619814, 
    -409.219771433257, 
    -547.152361392443, 
    388.266695958115, 
    244.502731420977, 
    368.008332909283, 
    660.806706623966, 
    370.102551318229, 
    537.276197563757, 
    446.717194287, 
    356.616614735807, 
    296.147245891953, 
    117.646995608513, 
    244.719400141035, 
    282.243533468726, 
    245.266593243211, 
    172.983336424108, 
    113.659337671714, 
    76.9067646220984, 
    100.020764205651, 
    44.9630689215159, 
    58.793600916462, 
    49.7442035482812, 
    43.4679406460828, 
    14.4616613829913, 
    41.7357350682607, 
    129.838930682132, 
    105.142879722099, 
    76.2971006075177, 
    122.282490680092, 
    159.036337458405, 
    206.110339432788, 
    293.244053971995, 
    301.378111152607, 
    333.305134063071, 
    416.918036487576, 
    429.753374029249, 
    566.070191027734, 
    618.770985405763, 
    647.728428070649, 
    686.487012796946, 
    946.223628737223, 
    1476.21561280663, 
    1590.78039516607, 
    1666.36154730136, 
    1409.2359019383, 
    1210.37636872874, 
    1168.97342892908, 
    882.1811024665, 
    1229.52139958878, 
    1.13387459204865, 
    1348.677910526, 
    -85.2539338254117, 
    -367.012049573533, 
    -163.84522470301, 
    149.675223304605, 
    405.777968168529, 
    582.67279099724, 
    413.968502642728, 
    463.344440481562, 
    -284.785340278172, 
    -304.87797179441, 
    -298.385892742025,
  
    -594.212571873511, 
    -544.750944583975, 
    -495.75030903747, 
    -444.136952813504, 
    -472.616422061558, 
    -480.885045140214, 
    -466.410364114691, 
    -491.764141804695, 
    -525.696857328512, 
    -520.053548934613, 
    -486.637934865238, 
    -552.053094665254, 
    -602.285427012343, 
    -673.497123402145, 
    -616.727980020994, 
    -491.391071870636, 
    -533.994142846316, 
    -23.1992412456777, 
    570.729430169849, 
    821.306133684626, 
    670.418095288593, 
    539.445182518357, 
    513.392227078873, 
    472.025681101597, 
    349.673352086665, 
    501.596449348988, 
    468.858324403325, 
    310.76239184543, 
    203.042757805362, 
    248.392729215633, 
    165.955394443714, 
    129.96537729714, 
    101.17100982196, 
    93.7005213430991, 
    44.9453683652377, 
    8.3478127591821, 
    31.1247329055117, 
    -10.3173938179342, 
    -1.92133849118186, 
    68.6421434251874, 
    25.7779304902798, 
    -43.5883724483925, 
    58.1773025302716, 
    181.716253870145, 
    167.577762922007, 
    244.97353076828, 
    277.501650332869, 
    308.761732872496, 
    438.671697883562, 
    543.412864193803, 
    506.934659404692, 
    553.967024697436, 
    643.260667858571, 
    657.96697541821, 
    783.27599024586, 
    1147.75369669369, 
    1666.61437931894, 
    1684.94567971908, 
    1386.49751083529, 
    1195.96585778455, 
    1055.62874065027, 
    1694.59667035794, 
    1710.60817796252, 
    1456.05882762127, 
    -10.1250552071126, 
    -283.960332913207, 
    -358.921820701437, 
    32.9016595346018, 
    243.547791012192, 
    546.032046558343, 
    150.041603094776, 
    580.74149711242, 
    27.8499547297775, 
    -239.574274522327, 
    -253.893046781704, 
    -270.246453557543,
  
    -746.002730118601, 
    -655.333342702765, 
    -617.45215807463, 
    -594.719213385331, 
    -564.76994524504, 
    -490.693557739258, 
    -501.324377361097, 
    -515.739515605726, 
    -539.958824157715, 
    -540.605010986328, 
    -528.904713680869, 
    -455.146671897487, 
    -490.162909859105, 
    -47.065276396904, 
    -55.654082398667, 
    742.649151551096, 
    280.5548111765, 
    38.3358132462719, 
    693.135076422441, 
    582.286392211914, 
    610.236457021613, 
    517.260599638286, 
    611.297836303711, 
    497.780514566521, 
    410.762183540746, 
    463.647856461374, 
    488.993668004086, 
    361.787082872892, 
    319.99027633667, 
    295.537562320107, 
    225.359699650814, 
    107.703618651942, 
    68.5944610896862, 
    50.1607074988516, 
    77.8580773504158, 
    27.652065129656, 
    -37.2334782951757, 
    -24.0913931570554, 
    -17.2362573523271, 
    -84.3328556763502, 
    -114.520487283406, 
    -116.237519264221, 
    69.7027043261043, 
    20.1802077293392, 
    81.644737067976, 
    212.265461369565, 
    158.134979549207, 
    263.629516601563, 
    299.975159494501, 
    414.032679507607, 
    456.690083553917, 
    525.482818201969, 
    522.828489203202, 
    609.090721531919, 
    886.676507648671, 
    1052.36001105057, 
    846.409101385824, 
    1565.39780064633, 
    1064.29564305356, 
    1595.37554690712, 
    1160.16508724815, 
    1490.75612278989, 
    2041.96448316072, 
    1749.88764311138, 
    556.93914072137, 
    -453.763794949176, 
    -163.968900680542, 
    142.360175986039, 
    246.352008116874, 
    517.643973501105, 
    294.17840114392, 
    641.776151155171, 
    -199.462251663209, 
    -241.779758553756, 
    -281.894914325914, 
    -287.480071419164,
  
    -846.866170714443, 
    -655.455321274573, 
    -593.233012209013, 
    -474.608990967206, 
    -488.388530641494, 
    -407.151154299199, 
    -370.664488857564, 
    -376.993948578701, 
    -360.727959012398, 
    -363.702193970376, 
    -319.923233702895, 
    -246.941552511388, 
    -147.144725199376, 
    -203.963641539399, 
    -407.228984405587, 
    -7.81818313344506, 
    689.342713436117, 
    572.638185456238, 
    629.770477602494, 
    1033.23496214727, 
    878.498415674635, 
    601.997862872458, 
    894.128676061001, 
    714.795584726707, 
    524.037249288527, 
    439.629138301495, 
    448.522335928205, 
    320.714612420435, 
    218.599765899334, 
    239.411371681752, 
    210.356784559977, 
    79.8118267603977, 
    30.4799012008462, 
    11.3326196173938, 
    -17.0866189214246, 
    -42.2680044347738, 
    -72.4702348340667, 
    -53.4866511229036, 
    -52.9166716309171, 
    -119.30404511865, 
    -127.791741137275, 
    -55.3119515091143, 
    55.5878302941533, 
    210.999532667547, 
    261.961377721618, 
    469.791676515962, 
    283.722394565185, 
    289.452037608369, 
    199.477470859302, 
    331.033465856401, 
    366.359654468225, 
    521.378257533605, 
    708.268542880308, 
    494.917584477989, 
    1014.03727786245, 
    1304.35681945186, 
    1275.83884194984, 
    1207.69559790599, 
    1559.64437418529, 
    1203.17112573023, 
    655.541360852972, 
    -262.601240899238, 
    -341.447027478214, 
    811.277141079795, 
    -581.363168963139, 
    524.960231400811, 
    189.213942203116, 
    358.856793705854, 
    412.505487465511, 
    497.747936663142, 
    432.266498813444, 
    180.717103721045, 
    -247.143183525573, 
    -296.212857206885, 
    -284.582547212368, 
    -469.621728407976,
  
    -971.549634397364, 
    -761.565436889717, 
    -518.968909004101, 
    -387.41263236017, 
    -382.784272718269, 
    -378.311969359805, 
    -305.86844092494, 
    -301.602050289995, 
    -280.207650708992, 
    -231.957946330943, 
    -129.794758573491, 
    -60.1930644606957, 
    273.870988087586, 
    389.806682932686, 
    -231.622525290706, 
    187.300331168589, 
    -245.079212393769, 
    337.792788698852, 
    1219.88537571172, 
    956.188148789012, 
    261.767732633053, 
    391.426470578183, 
    761.301501223915, 
    777.286329075043, 
    493.193072986495, 
    312.645090891292, 
    369.83170336545, 
    309.946217920318, 
    266.716157791462, 
    171.735969763453, 
    96.004005016698, 
    12.7388604909412, 
    -39.1900691238526, 
    -41.3245315023126, 
    -54.7623198558343, 
    -96.7478379103268, 
    -112.113672802189, 
    -96.9672791426553, 
    -50.1422831843975, 
    -43.488118976387, 
    -32.0094643157108, 
    -66.1504852918605, 
    -15.4978400996117, 
    169.812449628269, 
    549.676637382551, 
    307.227134593524, 
    425.902013058892, 
    414.605755258113, 
    314.012954617935, 
    280.878727783682, 
    314.590742989056, 
    398.633105484129, 
    782.427260805753, 
    1014.61567644416, 
    1176.16089781348, 
    1708.80146025757, 
    1509.42092340176, 
    1569.95509616899, 
    865.005692382681, 
    1256.44279032298, 
    -294.765298896796, 
    1012.60083139383, 
    854.319567476388, 
    1380.81035262873, 
    1623.65558119345, 
    940.932014807062, 
    240.867740671686, 
    803.00228574268, 
    636.448392135427, 
    500.365969543623, 
    505.454134207432, 
    -80.2367970424176, 
    -255.708808490971, 
    -354.987310595369, 
    -376.974396576407, 
    -587.818065480982,
  
    -1203.16666946326, 
    -976.527981697246, 
    -649.411338814696, 
    -405.03418430102, 
    -348.830867199187, 
    -327.700647467328, 
    -276.275188787787, 
    -250.684554032756, 
    -207.885823152634, 
    -203.502784444931, 
    -130.679392400274, 
    215.536769768692, 
    559.615714347643, 
    403.169278455609, 
    231.760076765255, 
    -8.44818787151796, 
    977.538336477246, 
    1150.38479507463, 
    1533.21670157165, 
    379.649434423934, 
    686.773067064279, 
    848.757252367455, 
    744.253433321519, 
    658.604449136526, 
    466.263279204673, 
    310.825949682768, 
    353.600589337835, 
    269.72303965057, 
    257.335953326935, 
    132.219050238674, 
    26.6219544434729, 
    -45.6251554029921, 
    -90.146366151423, 
    -56.4695331385531, 
    -80.2906741166839, 
    -111.185207176849, 
    -96.4691163583136, 
    -53.6374074929508, 
    -34.2203733010624, 
    30.132757339715, 
    88.7038127401512, 
    171.808120859965, 
    183.614704084024, 
    376.449310473606, 
    564.116843237456, 
    589.656969777414, 
    477.780285415563, 
    556.903543350545, 
    461.880842920113, 
    401.33134794075, 
    332.890383200309, 
    319.35808307353, 
    804.272699003663, 
    1204.91903860812, 
    1143.08596094352, 
    1500.31203582866, 
    1174.6698076135, 
    1504.62435050187, 
    890.681973815092, 
    354.829569723692, 
    1908.96448997849, 
    1627.07651580436, 
    2114.52344590686, 
    2094.74249479459, 
    1760.14860433854, 
    1102.72096088404, 
    900.15272197318, 
    501.754633212543, 
    179.05402046195, 
    146.351435033354, 
    100.866784919145, 
    -152.499088882199, 
    -252.404237486614, 
    -282.494834370202, 
    -370.389171719952, 
    -469.066038988205,
  
    -1611.64286488088, 
    -1141.3467852004, 
    -871.924097742506, 
    -532.223102855789, 
    -384.99537556596, 
    -311.585681095102, 
    -296.675765760535, 
    -266.092579456086, 
    -224.403807893179, 
    -196.598663451824, 
    -152.679176280372, 
    298.845471739904, 
    511.647721994366, 
    627.171526969749, 
    733.953582968721, 
    335.159746167908, 
    530.13359485895, 
    1682.79003593556, 
    1369.61233462412, 
    1460.73275030634, 
    1382.53845876115, 
    1083.21367400064, 
    900.069257558926, 
    642.552840152754, 
    557.651807855519, 
    501.55468985375, 
    443.610808723852, 
    337.725266899801, 
    247.609684071642, 
    150.417845863778, 
    61.3439724907226, 
    -24.3213996512084, 
    -65.7951905954323, 
    -67.7368251858206, 
    -104.579604934872, 
    -86.9524501200348, 
    -60.0626655265704, 
    -6.7803385410569, 
    19.5480055692544, 
    64.344475171601, 
    174.655560671817, 
    224.480016573814, 
    197.397972209456, 
    359.132865722075, 
    567.033866873782, 
    742.243474355872, 
    709.249641478262, 
    657.01157995995, 
    544.82697172261, 
    687.650382389016, 
    526.371908723975, 
    401.301126559131, 
    477.395501101539, 
    1037.29584421156, 
    1251.62478555677, 
    1575.21317256231, 
    1433.55325464333, 
    1637.23840275644, 
    1466.54858323255, 
    1874.64134327375, 
    1610.32236228678, 
    1558.07429757285, 
    671.110257711537, 
    812.932074364189, 
    1817.8274985182, 
    1053.74228438391, 
    1063.18045563394, 
    505.416189324017, 
    28.8722179364476, 
    89.0951051474449, 
    -191.657090883377, 
    -259.178120180581, 
    -252.475458568047, 
    -262.53913673922, 
    -263.551502898452, 
    -420.623614718103,
  
    -1789.02687906605, 
    -1480.3607293585, 
    -1016.06557389416, 
    -666.603964990357, 
    -430.661211532815, 
    -380.06345990684, 
    -310.623162422308, 
    -257.260733383367, 
    -226.1396849911, 
    -194.135756918724, 
    -130.92260706625, 
    -9.95450603254459, 
    185.282719730661, 
    301.77945493076, 
    1195.5172882849, 
    686.247723509989, 
    1099.08936869417, 
    787.139691778952, 
    1850.66317070665, 
    1388.73122907512, 
    1219.02629005629, 
    976.255105688215, 
    736.409365287686, 
    771.714932731125, 
    706.830242263777, 
    677.937988366686, 
    597.124433083869, 
    340.360144227509, 
    199.930438914198, 
    168.842260935272, 
    120.259644704863, 
    62.9736781435342, 
    -20.1613010756777, 
    -150.189165744376, 
    -18.5339261633811, 
    6.7701632790978, 
    -12.6114540204215, 
    139.866226637351, 
    90.3998308021577, 
    134.973160067705, 
    209.751169251702, 
    218.162846747864, 
    232.27159775438, 
    308.358244888459, 
    479.625278921437, 
    615.920283472421, 
    770.064786878972, 
    638.731708607774, 
    506.70408772194, 
    547.723955622177, 
    494.184512886995, 
    490.150542905323, 
    473.152704142778, 
    604.78351980895, 
    1052.79371939528, 
    1340.22726102105, 
    1210.49124620528, 
    1423.29658966235, 
    1778.02334874955, 
    1683.00844118603, 
    1852.42376474891, 
    1391.61756203239, 
    2054.10128367254, 
    790.234271315403, 
    1947.25909926189, 
    1083.21074239937, 
    794.997556483487, 
    403.364904939793, 
    386.853512105055, 
    -289.41337164252, 
    -375.367231794062, 
    -342.331181666085, 
    -260.773129361741, 
    -253.137120141161, 
    -284.553825207547, 
    -374.300028438932,
  
    -1945.78545882854, 
    -1664.82095381341, 
    -1290.52301283406, 
    -847.110106704216, 
    -513.385482664205, 
    -411.322031523052, 
    -360.68408303939, 
    -280.17285735503, 
    -233.228183154697, 
    -174.281872079727, 
    -210.276213768749, 
    -131.857944960555, 
    77.8856803284196, 
    822.567941074007, 
    903.734902573055, 
    644.920535626891, 
    1481.84492791701, 
    1788.1983496996, 
    1177.72859304669, 
    1154.00915390647, 
    1018.50771257458, 
    672.657356663751, 
    696.476776985945, 
    745.299268323123, 
    781.519781721399, 
    746.084410262669, 
    557.140511695376, 
    372.928654451786, 
    258.941471140436, 
    176.789129774087, 
    96.7839121065632, 
    53.3107246335381, 
    -38.8855371367098, 
    55.0678906721088, 
    -49.1641890516748, 
    -82.7436042456733, 
    46.0156986518515, 
    105.692102787876, 
    102.707225840142, 
    97.2606006207951, 
    137.166825227214, 
    204.35666732959, 
    260.017369448672, 
    307.134462371519, 
    382.742090393955, 
    511.359010788257, 
    833.617874743558, 
    871.099928348624, 
    563.047274095082, 
    569.902418540283, 
    749.266961844209, 
    685.074327441107, 
    871.370375894892, 
    975.569637678775, 
    1210.60912236708, 
    1437.11071931128, 
    1599.42469075066, 
    1412.93151195907, 
    1334.51244840376, 
    1216.87185053809, 
    1430.70302866288, 
    1254.76403731701, 
    1344.40184923195, 
    555.631260657223, 
    1195.19015911311, 
    321.182154972619, 
    11.2114740026715, 
    -326.256061842305, 
    -339.248701195966, 
    -375.718441996303, 
    -422.764237671921, 
    -394.233436780974, 
    -358.24406398504, 
    -311.218785801767, 
    -322.935276471488, 
    -455.790640046054,
  
    -2023.78228347966, 
    -1823.81358180201, 
    -1487.78491156259, 
    -985.96247997049, 
    -564.062797025231, 
    -439.692970946548, 
    -363.364166332386, 
    -280.88661151557, 
    -264.789370358458, 
    -282.292006269416, 
    -206.989840192463, 
    -159.304636052317, 
    0.581068660480788, 
    163.376427135705, 
    371.913781596458, 
    522.663495566782, 
    875.99170014145, 
    1300.27419064853, 
    1147.48452623801, 
    949.628202782232, 
    814.472341710481, 
    637.906652016976, 
    780.220826186366, 
    741.190680338313, 
    771.178674456521, 
    821.535642668755, 
    509.624031878531, 
    343.158281460854, 
    232.853265478255, 
    163.56735870686, 
    52.0488552563929, 
    -73.0641228749531, 
    -116.34085021601, 
    -18.5083461675008, 
    -64.9715160656083, 
    -76.7822206327379, 
    57.1054749216513, 
    131.493055761195, 
    173.378896527435, 
    87.1019993586604, 
    151.814905202937, 
    144.983007183264, 
    94.6641845767187, 
    232.119900082953, 
    328.475157632005, 
    495.513857001023, 
    879.094718625539, 
    1153.48566907518, 
    1057.28588856081, 
    822.041791396874, 
    900.183540839768, 
    918.069312049721, 
    855.708413990189, 
    1071.87676802034, 
    1139.67965983597, 
    1354.09223309182, 
    1534.01393778461, 
    1650.23781403715, 
    1090.46179007843, 
    1376.89989303128, 
    1513.90697779127, 
    671.951665316586, 
    1457.28702887762, 
    1140.5978653877, 
    -118.913752364701, 
    -335.886622207826, 
    -114.541111479408, 
    408.565448450756, 
    310.449693143698, 
    -94.0047174749577, 
    -200.289580777671, 
    -206.154594498278, 
    -238.99376543265, 
    -243.02389974263, 
    -275.64627437442, 
    -322.1150713597,
  
    -2103.3155948515, 
    -1949.38589041818, 
    -1666.07602313171, 
    -1239.94000213384, 
    -749.927712657285, 
    -380.172740201533, 
    -308.181962751194, 
    -320.868107551157, 
    -313.298585522215, 
    -266.225705248243, 
    -318.290922226858, 
    -356.701568787203, 
    -160.199857203715, 
    310.819853347998, 
    417.796067954451, 
    570.881670858933, 
    665.951244589195, 
    776.395693506664, 
    707.74600834008, 
    765.462486121848, 
    651.646086851933, 
    561.604531214458, 
    708.151252387753, 
    680.386389677895, 
    654.366071233289, 
    571.508961488523, 
    371.668007653076, 
    315.799154604135, 
    278.457924538471, 
    164.602011412549, 
    70.3144347227164, 
    -43.7959824804495, 
    -144.660031095464, 
    -58.8091336733025, 
    -91.5506393906789, 
    -13.2545724173509, 
    41.4180403722228, 
    108.109840386658, 
    169.089018656185, 
    172.929502863099, 
    174.211155796371, 
    152.17686819523, 
    124.494167375939, 
    147.293880906912, 
    275.549333948305, 
    601.112536269103, 
    855.527202960759, 
    992.219325775794, 
    867.897983768878, 
    804.0465274311, 
    1049.03015827038, 
    1058.33867060885, 
    964.273518202421, 
    1423.96860055614, 
    1506.38472049794, 
    1153.31007294692, 
    1881.30061822188, 
    2145.91047800028, 
    1584.42769580939, 
    742.29598770054, 
    1222.37769446634, 
    20.1675171035037, 
    1278.20503528761, 
    1012.16331100036, 
    -272.080478856175, 
    441.767511698863, 
    299.701729551269, 
    136.785158052691, 
    256.353480229061, 
    -181.614274782138, 
    -228.071485745813, 
    -241.323742248177, 
    -253.976599683687, 
    -253.406795732385, 
    -254.075100180016, 
    -357.057773406402,
  
    -2165.34945798321, 
    -2049.73871774022, 
    -1777.27532232782, 
    -1324.35465323351, 
    -867.049110489489, 
    -354.200272729922, 
    -293.003040130034, 
    -299.822773001095, 
    -247.747864974172, 
    -223.861479738926, 
    -192.779951283538, 
    -287.829655347184, 
    20.9800124496101, 
    220.173360531975, 
    99.2917163855287, 
    182.378237857792, 
    315.992727311698, 
    460.588516222533, 
    484.458528174796, 
    497.402968198426, 
    553.362651974462, 
    676.030437405406, 
    634.171655541703, 
    547.397012699891, 
    498.813022634883, 
    367.3903851995, 
    225.823093717603, 
    231.50834486172, 
    209.523416884401, 
    177.359952834793, 
    118.049733259109, 
    0.945912824032069, 
    -123.914423801597, 
    -104.390110588287, 
    -27.7747263417131, 
    -9.28324343267445, 
    7.61740910579704, 
    -39.8032659007224, 
    48.835236330448, 
    94.2061285849778, 
    152.737862812311, 
    138.128201799723, 
    157.161980454892, 
    120.936379417727, 
    315.381259023278, 
    777.829054222662, 
    674.574206165341, 
    794.484657287597, 
    684.072456675977, 
    983.045347463649, 
    1240.86671517811, 
    1128.58557788469, 
    918.356785696274, 
    1612.01461568151, 
    1360.98831718419, 
    1762.68155917075, 
    1934.54893105775, 
    1811.49847729932, 
    1773.98137525535, 
    688.15821715354, 
    1461.68418316985, 
    1248.39027808039, 
    376.576893980554, 
    309.195147028424, 
    703.609463354263, 
    842.698802798475, 
    472.929830997543, 
    27.1516045245166, 
    -104.281339771404, 
    -199.823249731459, 
    -306.668656412193, 
    -322.36093974781, 
    -255.788843268109, 
    -256.007186377035, 
    -262.908270772867, 
    -376.57775729394,
  
    -2180.35901111291, 
    -2058.27014431841, 
    -1775.41798182164, 
    -1116.44831189436, 
    -634.196946899141, 
    -417.080525239132, 
    -318.623618131256, 
    -276.896543855229, 
    -186.818966176715, 
    -186.153864637334, 
    -194.938682966243, 
    -197.960014104042, 
    14.1367075180245, 
    42.56986832325, 
    -3.2713918027463, 
    -74.5708094326642, 
    303.588835053058, 
    438.368874497538, 
    344.701644594165, 
    381.665694481315, 
    449.124616748946, 
    562.895974102639, 
    451.925863225408, 
    420.898550133955, 
    409.80788938943, 
    298.956398262288, 
    234.820699824196, 
    254.107172616786, 
    227.920424643983, 
    197.679800178809, 
    72.351860558999, 
    -23.0686332441255, 
    -116.860569517129, 
    -182.060407397196, 
    -47.8119345683131, 
    -25.9278356687221, 
    -18.3663366751337, 
    51.3756185325501, 
    26.6282099831145, 
    14.8419516209382, 
    -17.7673961335323, 
    38.9904779899281, 
    44.7565404992341, 
    164.086529989126, 
    397.946602367477, 
    527.111475492784, 
    420.37650312742, 
    673.46920743902, 
    932.187488953184, 
    1173.19931124253, 
    1307.84514777684, 
    1292.97715687511, 
    1331.31702295797, 
    1674.79194736801, 
    1654.79951365985, 
    2114.61573909405, 
    1967.38433038212, 
    1890.85328850313, 
    1598.52536777954, 
    518.210159010774, 
    187.539078817141, 
    1327.95503457847, 
    812.285014623463, 
    -106.793885676919, 
    497.584438080479, 
    730.870181939118, 
    386.651882171645, 
    376.119465890953, 
    -17.9124088910458, 
    -194.444099212683, 
    -301.413391023574, 
    -202.671166773472, 
    -246.320677922795, 
    -263.68745743601, 
    -255.340687028772, 
    -306.651770951632,
  
    -2202.69079309615, 
    -2029.69510046605, 
    -1570.34760556963, 
    -903.620491788206, 
    -651.67046797903, 
    -577.461472335082, 
    -475.689799185966, 
    -336.894155448923, 
    -186.114302743056, 
    -128.798963343843, 
    -178.193308859097, 
    -281.688430850208, 
    -14.420464014953, 
    48.8236599914643, 
    177.997332630612, 
    297.110419197556, 
    363.265599676901, 
    392.123255256578, 
    374.467734235398, 
    357.562551154535, 
    349.404056903627, 
    504.357259842209, 
    443.652987506862, 
    397.253404051299, 
    380.013952693106, 
    316.057112015642, 
    184.757820870548, 
    153.502878449665, 
    142.881286864583, 
    101.963678350373, 
    52.1076125249615, 
    21.7513869954117, 
    -138.716844237267, 
    -303.468883766439, 
    -79.2471253495459, 
    -30.5654820733753, 
    -66.1793362696526, 
    -83.8279564020224, 
    -34.5514869545778, 
    -33.1188168312116, 
    -88.902761332266, 
    -53.5497325046061, 
    158.378381562531, 
    215.773679733277, 
    127.603204075721, 
    559.24668960315, 
    651.987902300618, 
    700.189398745274, 
    835.329863809924, 
    1185.37438264272, 
    1150.48424131045, 
    1453.27684752324, 
    1246.60302763424, 
    1791.94634556958, 
    1979.44179954401, 
    1950.8578814499, 
    1673.69428400976, 
    1815.16271832542, 
    1224.95637934257, 
    575.710524239675, 
    340.197603320243, 
    772.92325869921, 
    1294.30115169853, 
    771.233730628001, 
    710.496015362888, 
    481.691730225883, 
    -37.9806164680735, 
    -13.8464572421709, 
    -171.225253974474, 
    -261.332047636537, 
    -219.862207961642, 
    -207.483444647453, 
    -238.522488870652, 
    -256.324912431125, 
    -255.447367812324, 
    -262.417451038339,
  
    -2200.83328992068, 
    -2053.71045249948, 
    -1449.89971758083, 
    -969.48091075081, 
    -655.949930991996, 
    -700.545485083227, 
    -652.570897144009, 
    -581.557467325006, 
    -391.758307680175, 
    -204.502747312509, 
    -337.307414367782, 
    -417.57518263387, 
    -102.430272003839, 
    23.7457414354232, 
    152.227516966999, 
    304.871008579301, 
    349.068916564293, 
    283.68763915315, 
    361.464465971092, 
    401.535951800203, 
    464.813461047405, 
    486.997526657941, 
    437.94686847785, 
    399.072588041675, 
    345.62022608365, 
    337.008955277361, 
    244.133816688085, 
    154.333632177629, 
    78.1036647228502, 
    93.5517135867878, 
    58.6868053598604, 
    20.0390427258084, 
    -77.4167477617349, 
    -258.264453986189, 
    -100.641786007171, 
    -83.3909046999693, 
    -128.145574313397, 
    -136.772941230527, 
    -150.205379289583, 
    -115.933661284667, 
    -111.905313250466, 
    -88.1336206434029, 
    216.551175214673, 
    247.916178492921, 
    229.378074861721, 
    398.484548293198, 
    753.265779168453, 
    627.535317441249, 
    561.100375449933, 
    780.983324552834, 
    1208.28314953983, 
    1181.19042493727, 
    1278.16429978869, 
    1727.02453861044, 
    1825.91958182442, 
    1992.96159822436, 
    1816.12746924115, 
    1997.42543557777, 
    1842.19079331829, 
    1112.87048613238, 
    1783.03023555539, 
    1398.89508355665, 
    176.469551423345, 
    852.788603557314, 
    738.699896373509, 
    -65.586197699863, 
    -328.91231893986, 
    -359.128282258653, 
    -103.371631600949, 
    -144.71966949796, 
    -194.165727329148, 
    -196.409777524891, 
    -199.395623727182, 
    -286.905601091375, 
    -293.2546673056, 
    -278.60635333686,
  
    -2180.47908524089, 
    -2063.91038649881, 
    -1729.5092844349, 
    -1100.37124197213, 
    -649.384470940705, 
    -438.83400413197, 
    -604.498825628573, 
    -644.327571856081, 
    -741.847952275634, 
    -749.361830204092, 
    -711.984812011377, 
    -349.185611235735, 
    -70.4761397016272, 
    55.8481818361481, 
    62.8948240568493, 
    249.628612889955, 
    245.375755083654, 
    221.565399896124, 
    401.13328638536, 
    419.449543836536, 
    431.832943505162, 
    501.351527966951, 
    445.143663908306, 
    412.347887801697, 
    346.758902563627, 
    354.766676472389, 
    281.229605556202, 
    198.72266503491, 
    159.913706718607, 
    104.597610511011, 
    39.0169758719262, 
    37.6033038863409, 
    -59.3200748118953, 
    -163.89528107296, 
    -139.738859057026, 
    -120.604329586563, 
    -170.028645149137, 
    -166.23815598867, 
    -175.453650919881, 
    -203.180799379594, 
    -41.4751681373723, 
    -55.7283377444492, 
    62.863653132725, 
    58.6979392148876, 
    -37.6154900189879, 
    355.991094685352, 
    772.878975324642, 
    496.635256422323, 
    299.70406048936, 
    524.73967590845, 
    990.208869754667, 
    815.674191055211, 
    1037.02443231154, 
    1489.09764799693, 
    1569.96135816755, 
    2083.86521756129, 
    1796.15689285124, 
    1549.49195496152, 
    1115.07752404635, 
    1708.70219939126, 
    1750.60231566563, 
    1479.61781599807, 
    497.726460908586, 
    -49.3851008196332, 
    110.345900417046, 
    845.315759878812, 
    838.575950297904, 
    46.2948742051659, 
    -312.916203254281, 
    -323.359122563584, 
    -366.119608230848, 
    -419.788486903619, 
    -363.939216724836, 
    -389.860282453685, 
    -356.864954770078, 
    -346.134432054714,
  
    -2155.92419935955, 
    -2046.99928743335, 
    -1886.83335505675, 
    -1466.96730181618, 
    -622.443630957523, 
    -423.295896792866, 
    -330.840162736438, 
    -389.067571253418, 
    -524.050514627009, 
    -688.300373320883, 
    -860.895256871205, 
    -390.125334484448, 
    -73.6002514108696, 
    -0.0193961415885698, 
    168.920977128982, 
    337.455960708397, 
    178.911351145181, 
    53.897756860077, 
    347.68496435834, 
    425.968928816604, 
    490.780634915308, 
    507.482119296458, 
    348.03373531585, 
    396.93212763326, 
    351.190681017526, 
    325.40977630957, 
    213.89334938374, 
    200.139024975852, 
    196.121607313765, 
    110.458186712404, 
    90.001177494096, 
    43.980462030227, 
    -30.4211546523041, 
    -56.7264338191117, 
    -61.0345540276301, 
    -126.667538590554, 
    -161.44704077145, 
    -179.950858238964, 
    -169.039298088527, 
    -130.35828568073, 
    129.538699111641, 
    50.6481944080966, 
    -101.609387589996, 
    -67.4943473523301, 
    34.8858221484997, 
    264.769282506536, 
    670.416852320963, 
    166.276554635225, 
    524.019761080174, 
    1113.17772232859, 
    1164.02765135215, 
    816.875218330544, 
    825.99240455756, 
    1473.10773436407, 
    1814.333393161, 
    1878.10579208938, 
    1884.08312055325, 
    1576.64809052915, 
    1817.70732767718, 
    1498.97792306112, 
    1189.00293628313, 
    332.248882716616, 
    592.194333613653, 
    -84.7180286612538, 
    655.635504416089, 
    649.794365732301, 
    370.925762338839, 
    108.142810731825, 
    100.882016439854, 
    -165.13118797721, 
    -275.78691319362, 
    -298.179507149827, 
    -249.26750940278, 
    -252.118518842161, 
    -296.636093618087, 
    -298.210120360234,
  
    -2136.89420304079, 
    -1998.67952173795, 
    -1794.29047744939, 
    -1138.29368261527, 
    -385.782996042044, 
    -366.042017929231, 
    -378.131436013695, 
    -277.189188706247, 
    -276.188354808298, 
    -283.081576408222, 
    -697.597856912474, 
    -571.607610862708, 
    -25.9949688169207, 
    71.6634131172055, 
    149.087289395816, 
    361.009920887023, 
    241.863295402398, 
    121.557694618806, 
    238.704457501949, 
    339.560510868187, 
    429.714982860432, 
    473.976005067217, 
    321.347796774391, 
    321.931245549663, 
    327.634463260048, 
    304.790904323838, 
    213.881858114432, 
    154.258716100541, 
    115.29958045229, 
    54.2424037218891, 
    55.8676401241897, 
    37.529269077743, 
    2.69196665760915, 
    -27.2569167322969, 
    -79.9444199921973, 
    -158.410887142579, 
    -177.848794307046, 
    -169.736350594549, 
    -145.417072657107, 
    -102.899801750866, 
    -8.28343940909221, 
    43.4906405975404, 
    -43.629790594704, 
    -77.4666823561219, 
    -43.1119641974682, 
    187.737865131888, 
    262.207444307385, 
    108.257514689831, 
    530.194503690202, 
    1001.10385400958, 
    1078.07956171837, 
    644.654836092923, 
    879.81928276242, 
    1453.65748252741, 
    1628.62383939224, 
    1678.22556821816, 
    1799.88439796166, 
    1767.38742362745, 
    1508.0504726568, 
    1268.6431230671, 
    920.512978984155, 
    1241.17461442253, 
    780.976300084702, 
    352.324112794969, 
    1017.66604814177, 
    887.086602820795, 
    693.366909919907, 
    428.16156991786, 
    387.796451923158, 
    -43.1060434944307, 
    -145.387265014222, 
    -172.765044676897, 
    -200.760280265253, 
    -203.73652383862, 
    -232.452664421227, 
    -271.426373997567,
  
    -2211.41779924587, 
    -1938.75389861206, 
    -1455.13970157841, 
    -572.275736724407, 
    -406.82123109448, 
    -395.094517898987, 
    -376.470691958574, 
    -342.601219950438, 
    -288.43981515814, 
    -152.13046942366, 
    -350.786529609364, 
    -555.693122389603, 
    -164.536226877039, 
    227.282547153522, 
    76.4381926842, 
    353.981681708393, 
    224.448014745252, 
    149.937925419909, 
    185.367049773623, 
    264.069068325594, 
    391.481390872969, 
    382.949499593736, 
    383.133342452439, 
    400.245082547657, 
    312.588338303005, 
    240.443639665541, 
    209.552355002716, 
    146.547851871135, 
    177.694932410058, 
    191.397038599679, 
    66.0745562839614, 
    30.1967093322473, 
    17.0861820018571, 
    -25.6782364925372, 
    -102.641237492791, 
    -129.93965312962, 
    -137.178414377894, 
    -144.476428801909, 
    -89.2459704814537, 
    -72.1341166223948, 
    -98.1447306127857, 
    -67.4112487731026, 
    -58.3726805791609, 
    8.24141975132699, 
    63.0131255755375, 
    263.339604380951, 
    316.206085952638, 
    111.953999458476, 
    494.994132342025, 
    828.639969119834, 
    771.951281625505, 
    740.051637579053, 
    1123.97526907414, 
    1243.52241471687, 
    1457.57506941468, 
    1510.84000561619, 
    1446.94528304181, 
    1606.84386716631, 
    1495.83967720194, 
    1468.91146472961, 
    1113.67458178615, 
    240.805139330173, 
    395.825438235667, 
    500.999642289892, 
    686.413738891495, 
    1222.48520438269, 
    227.495050491166, 
    955.892539636286, 
    442.081719397431, 
    -54.4957391031665, 
    -165.089389422974, 
    -188.534162066418, 
    -244.760768080879, 
    -231.149673812199, 
    -273.141074066333, 
    -331.90351339684,
  
    -2065.35657500366, 
    -1776.82241764902, 
    -677.686365133968, 
    -469.971555588094, 
    -479.334462480877, 
    -483.779356402219, 
    -453.857910015282, 
    -423.748358988148, 
    -358.461440783733, 
    -208.522038033668, 
    -140.013935441533, 
    -336.034984216979, 
    -156.010856551526, 
    -3.18785507441785, 
    193.872155992074, 
    326.630434525372, 
    66.0682818011238, 
    159.357590986126, 
    163.556632630369, 
    268.190894899016, 
    406.487380866108, 
    468.211177415837, 
    490.426445613917, 
    431.800428533607, 
    303.761887681711, 
    234.733440330822, 
    140.408850378312, 
    165.353422570737, 
    273.061984041904, 
    293.094624437116, 
    161.382187007122, 
    70.3990697396164, 
    52.250426878721, 
    -4.20739397089523, 
    -126.021618371047, 
    -132.244014963191, 
    -116.798047547378, 
    -95.4089778289278, 
    -86.2332362947109, 
    -78.3346997054934, 
    -63.4611004373394, 
    -47.5057555798855, 
    55.2841320898631, 
    -23.163215096827, 
    -1.42829508276895, 
    89.7515443447329, 
    291.612068381316, 
    357.640793495991, 
    521.127139750412, 
    786.080950951655, 
    475.468806972695, 
    672.43599324157, 
    915.805118360019, 
    1210.6751683012, 
    1434.2324068896, 
    1551.29165234197, 
    1521.99660381731, 
    1471.40814962526, 
    1533.91442845463, 
    1520.59315671846, 
    1436.20499402225, 
    1184.59230572912, 
    1021.35713891246, 
    923.727482401648, 
    579.706465931507, 
    434.20012717765, 
    2.22718926186129, 
    32.587657339628, 
    -194.031711445945, 
    -147.719466263614, 
    -152.960954755846, 
    -205.733434730521, 
    -239.196241541113, 
    -266.350792396776, 
    -276.026307480867, 
    -273.559281531801,
  
    -2111.80135452253, 
    -1581.50265128722, 
    -592.309491404228, 
    -565.822331709398, 
    -559.197528433293, 
    -567.289305128416, 
    -517.653068123847, 
    -518.813582391515, 
    -499.102194142102, 
    -378.324367360868, 
    -157.568376075515, 
    -356.24707617338, 
    -101.536068539337, 
    -7.13024460942492, 
    153.767326504489, 
    178.753336914975, 
    280.912307239461, 
    337.469319961907, 
    188.760851301513, 
    358.90147730538, 
    334.849052202795, 
    382.713426989377, 
    556.959217306483, 
    534.162522618208, 
    428.229850380312, 
    321.026557875374, 
    246.736715474828, 
    307.589020522952, 
    299.728109562651, 
    260.657148728578, 
    166.728495838126, 
    110.571743147104, 
    61.1016791900084, 
    -12.7650181795601, 
    -191.765516063267, 
    -118.938118227652, 
    -122.392013331944, 
    -50.9165407679514, 
    -50.7719686738855, 
    -45.9264016332977, 
    -36.9149328912098, 
    -139.003535808935, 
    -28.4185347145913, 
    -47.2419231244994, 
    -47.6014838005098, 
    163.946604068712, 
    450.709277243792, 
    475.145656261038, 
    402.363573354142, 
    410.737806638436, 
    385.79871598657, 
    536.860564104787, 
    851.924878717402, 
    1001.91159342972, 
    1119.22125452603, 
    1350.64600878948, 
    1466.16063209183, 
    1008.19100659958, 
    1289.60449071801, 
    1687.03005422697, 
    1698.6094103874, 
    1649.97740988394, 
    968.555392881525, 
    707.838196937065, 
    631.613575378979, 
    480.299594422069, 
    756.517842394244, 
    957.2839564615, 
    9.85369958535791, 
    -268.424895360249, 
    -235.091731993109, 
    -233.395891223749, 
    -299.307175477167, 
    -231.127709268055, 
    -242.337750089929, 
    -304.836555322902,
  
    -2179.75245200026, 
    -1527.17341007177, 
    -693.530680589154, 
    -677.690123144751, 
    -657.223130818845, 
    -629.967502700789, 
    -585.229425863884, 
    -552.117259231688, 
    -596.946277255307, 
    -603.757409603039, 
    -491.135614025636, 
    -514.959440353068, 
    -155.847855594631, 
    3.11219056549723, 
    78.8367592778476, 
    104.463709534351, 
    257.596890230595, 
    326.131119410911, 
    271.859755388966, 
    405.789939649695, 
    374.755217826647, 
    528.227008806767, 
    670.477693641039, 
    613.48771058325, 
    479.072214376486, 
    357.178319360748, 
    300.34700288591, 
    369.334636636971, 
    293.741968682472, 
    178.395095776069, 
    150.322375627541, 
    131.687876773975, 
    72.9764484440758, 
    -33.0310216310447, 
    -202.022645014798, 
    -124.39851581236, 
    -136.058407105364, 
    -98.8480887578561, 
    -97.4379493835128, 
    -101.297125929548, 
    -15.9852761026182, 
    -12.2511925963812, 
    -21.8187641438023, 
    -94.5891343572781, 
    39.3187287729519, 
    353.035763820636, 
    432.864687203027, 
    539.610340848881, 
    450.986482511309, 
    363.400185024352, 
    389.638995325446, 
    439.902814995402, 
    557.80479625091, 
    612.342069465661, 
    955.386850619768, 
    1234.54740095833, 
    1113.51298193168, 
    1198.38130321268, 
    1202.85594735994, 
    1364.20279366385, 
    1352.39918970874, 
    1002.66878985397, 
    813.467199848854, 
    1166.4113264949, 
    1456.73090452257, 
    963.054791799706, 
    343.566253946181, 
    562.76868390876, 
    137.314656286735, 
    177.124143994337, 
    -183.052361527856, 
    -198.391019020209, 
    -169.660394228586, 
    -210.022562372992, 
    -225.611264236296, 
    -402.533418033852,
  
    -2247.27028291196, 
    -1583.30900378938, 
    -851.591013114905, 
    -755.201975310904, 
    -703.302779792538, 
    -642.944580556563, 
    -623.559665786726, 
    -621.948821679743, 
    -660.012693783204, 
    -710.300371048298, 
    -782.830360147748, 
    -688.463677349709, 
    -102.827791204377, 
    -3.27704165096856, 
    47.5599633141537, 
    140.515364867978, 
    189.150340457245, 
    244.225375578089, 
    206.405992067942, 
    494.295485856419, 
    582.535712358533, 
    614.887783627227, 
    647.721790292361, 
    657.917014067544, 
    523.115379478737, 
    379.012372840291, 
    348.698252435493, 
    416.499344918656, 
    258.447858201696, 
    115.84423148592, 
    173.134796112676, 
    131.158101155536, 
    68.6210361584291, 
    -82.4972280970083, 
    -120.123252971174, 
    -111.094600589919, 
    -131.248547382077, 
    -121.440820281743, 
    -84.9859663492362, 
    -114.098828655341, 
    -99.5118684747326, 
    -93.1662727518298, 
    -191.49832717195, 
    -196.73697434027, 
    -57.4619000799048, 
    190.600170506075, 
    382.579643651058, 
    473.965219375935, 
    543.177241702363, 
    572.294850920778, 
    605.157894702668, 
    499.326417600455, 
    506.758384644785, 
    409.721317047769, 
    671.38051331831, 
    998.306511489166, 
    984.015477350275, 
    771.855668028421, 
    900.83748449003, 
    979.013206507566, 
    1255.50161965297, 
    815.85593962803, 
    1014.7043536999, 
    1555.67494886853, 
    876.617178298581, 
    1200.05721165913, 
    740.38562417538, 
    581.402118524811, 
    276.338229586267, 
    257.243494601951, 
    -152.46378639751, 
    -164.21199135177, 
    -210.0775943, 
    -211.915795410601, 
    -211.117755434948, 
    -313.148394925329,
  
    -2259.70886086937, 
    -1842.85755325779, 
    -1056.1645660144, 
    -803.557179988164, 
    -737.672263654855, 
    -686.589854890795, 
    -644.972457484197, 
    -630.344661802354, 
    -696.373624299702, 
    -754.968976284596, 
    -806.802819930159, 
    -527.66430885768, 
    -102.831578559598, 
    1.84802969846306, 
    1.74380039177536, 
    235.705879897047, 
    174.26799510815, 
    251.80043602417, 
    335.618584435305, 
    484.466067571524, 
    500.100097895468, 
    470.584562619881, 
    511.968336440679, 
    461.691237211491, 
    480.997039735116, 
    401.266300227049, 
    396.464553072632, 
    333.318388756283, 
    155.05308021383, 
    166.984178980948, 
    158.614638526121, 
    79.7821655679249, 
    -35.6451787148999, 
    -115.1972951857, 
    -110.497508951425, 
    -133.260885870871, 
    -133.997083890345, 
    -138.640179654386, 
    -141.773622104863, 
    -95.9790077711405, 
    -200.725428934728, 
    -177.527195517187, 
    -163.769643042415, 
    -137.765398416379, 
    -113.619305800749, 
    105.248540501312, 
    215.248358315342, 
    414.933467702664, 
    619.518490294728, 
    590.612745654542, 
    545.706826999232, 
    480.184057891435, 
    643.484632084114, 
    690.419392371099, 
    770.415488940472, 
    828.874181706855, 
    855.980757804097, 
    913.537974068185, 
    995.867957504979, 
    1352.12875781428, 
    1272.90640674005, 
    1149.3168106848, 
    1363.82231343474, 
    1558.3327285066, 
    1234.94789228622, 
    947.001989067738, 
    583.146869578258, 
    104.455097432637, 
    -125.859225099058, 
    240.476212961815, 
    -139.477781953631, 
    -215.627962669894, 
    -217.180597320249, 
    -251.714147642506, 
    -268.339031794037, 
    -275.91311424657,
  
    -2241.84539186621, 
    -1922.83363682319, 
    -1305.77318443991, 
    -775.655602902608, 
    -418.940517493885, 
    -317.716048634732, 
    -530.986292494101, 
    -676.340110727547, 
    -737.207844374296, 
    -758.954282070728, 
    -832.47850480886, 
    -559.878123032422, 
    -156.623840815811, 
    -6.7596271259658, 
    119.400227945038, 
    102.352621596975, 
    102.249843400374, 
    283.896625653361, 
    444.002198683855, 
    520.152608557483, 
    476.412861741805, 
    396.869970302432, 
    326.15504971597, 
    313.389108877833, 
    393.26148495989, 
    448.115299835716, 
    363.73785387148, 
    293.935033198032, 
    130.686745643616, 
    114.672511663575, 
    125.751152977297, 
    46.0165735495183, 
    -79.5553426667801, 
    -107.183069181068, 
    -136.489986218904, 
    -157.39974030028, 
    -158.68299919547, 
    -150.430320047718, 
    -122.658518606444, 
    -69.2584982911523, 
    -106.754997646421, 
    -59.5228298391211, 
    -61.7921846015715, 
    -78.8723210690398, 
    -38.4673629896365, 
    133.043331544585, 
    213.178846412651, 
    391.516257915092, 
    580.169509605755, 
    430.335380942929, 
    504.341519085584, 
    374.72352002476, 
    580.202045444948, 
    786.604986919136, 
    769.28010090041, 
    877.017315043317, 
    918.067534452059, 
    850.844640152992, 
    800.269045437842, 
    765.505884048787, 
    996.996295403528, 
    1169.04996528925, 
    1263.45085272196, 
    1303.05323080679, 
    847.160409873963, 
    305.700736202821, 
    424.823914710502, 
    240.184993089236, 
    -201.302951445373, 
    -193.704892986168, 
    -188.021388783305, 
    -255.48638630661, 
    -286.888877390214, 
    -299.7344196059, 
    -298.826346419827, 
    -299.694674531396,
  
    -2230.45114101568, 
    -2164.57618926968, 
    -1704.00540434527, 
    -963.784400196653, 
    -560.094707424937, 
    -326.418264972136, 
    -446.871469093995, 
    -463.938504841665, 
    -705.509915675452, 
    -753.630387975815, 
    -796.202511965761, 
    -420.230666037768, 
    -198.27578607839, 
    -55.4214073922863, 
    -221.542091183811, 
    16.3659481180633, 
    187.9049543061, 
    292.638145305808, 
    450.97037379659, 
    397.680835843488, 
    288.96955323086, 
    254.652184626293, 
    334.766162756978, 
    301.699260737302, 
    309.46417521256, 
    447.309089105315, 
    345.206393905078, 
    275.8109007939, 
    129.650452755867, 
    15.08072540995, 
    83.3796849309541, 
    37.0132770132497, 
    -120.676918631038, 
    -88.7508215439683, 
    -151.642689917416, 
    -155.27729391758, 
    -112.61548067928, 
    -117.828685695353, 
    -105.649036048641, 
    -61.4920234146202, 
    -79.9214676406336, 
    36.5347513698652, 
    126.611843636696, 
    94.9206034862196, 
    122.479610998447, 
    211.235866347995, 
    192.925968204339, 
    353.666549682617, 
    394.428256275137, 
    281.432979938297, 
    407.972438927593, 
    409.798844366298, 
    595.605651052378, 
    895.650187698482, 
    942.330175094349, 
    1102.1582098317, 
    831.939598655913, 
    1127.3830092239, 
    823.2497320912, 
    649.057623304698, 
    1055.01288525281, 
    1180.94031233324, 
    1541.57855875629, 
    1517.97635648071, 
    917.204163486175, 
    928.562512798248, 
    -86.3399059620251, 
    -328.141804194262, 
    -256.700441037949, 
    -206.016915422796, 
    -280.020204781149, 
    -338.800892141071, 
    -361.069677859112, 
    -314.771796979402, 
    -271.243946216407, 
    -208.48919670045,
  
    -2211.78012676175, 
    -2191.58434942401, 
    -1785.7442736994, 
    -1001.021441418, 
    -433.203738094042, 
    -305.447157049232, 
    -244.995249659588, 
    -420.024059658756, 
    -628.952746247123, 
    -806.044024203687, 
    -698.3559857974, 
    -435.941152327005, 
    -195.39898460149, 
    -46.5513604854018, 
    66.1165585993143, 
    169.840521463218, 
    240.410581103895, 
    263.813337849343, 
    422.701433542725, 
    540.185764052165, 
    576.75845598347, 
    544.089490217699, 
    423.980027706065, 
    381.391899066167, 
    500.705020391926, 
    448.233777724348, 
    378.256685425693, 
    321.876777153398, 
    198.443657083716, 
    204.551753769265, 
    128.483438781234, 
    -15.4782488227286, 
    -136.918456270872, 
    -94.5413402822227, 
    -172.813598201365, 
    -180.075673980115, 
    -158.966916087494, 
    -161.438109524974, 
    -124.333487069621, 
    -61.4766303966985, 
    -29.64342207831, 
    47.5001464381345, 
    118.111227120958, 
    104.267587049811, 
    102.282105624209, 
    197.280806914154, 
    120.079447524144, 
    146.314382695133, 
    176.156511889858, 
    163.330899587804, 
    322.104046948679, 
    421.234599131619, 
    600.817564807307, 
    709.784956501683, 
    815.123357578461, 
    1097.7215157025, 
    847.603322378332, 
    1272.27669927548, 
    1283.39346844886, 
    1283.22443149819, 
    881.878573085523, 
    1131.41496746752, 
    1525.07522429224, 
    1065.84414570328, 
    1017.62083582007, 
    253.464526113463, 
    -93.6812083670322, 
    80.6084682148488, 
    -29.8323455246655, 
    62.2724990567057, 
    30.5902993804584, 
    -262.453880393358, 
    -324.95237745176, 
    -261.560052948595, 
    -209.319215580169, 
    -193.414416690156,
  
    -2180.25489453426, 
    -2133.83683604276, 
    -1343.94542454017, 
    -580.312760715116, 
    -342.738302455103, 
    -239.79324165891, 
    -193.882169702151, 
    -353.661117156432, 
    -623.06314255222, 
    -855.356810224818, 
    -692.614686395662, 
    -216.440216606968, 
    -193.814234839308, 
    55.8967354091963, 
    340.255908054051, 
    274.498757453148, 
    264.069895202881, 
    353.781864871106, 
    448.179210842261, 
    396.333445558625, 
    552.123931355065, 
    514.881611455594, 
    393.619855451423, 
    309.308703756816, 
    342.44874770537, 
    328.678260072746, 
    353.43604691218, 
    331.919479357301, 
    245.200858055277, 
    185.886728261111, 
    67.7405661618162, 
    -34.0290391517253, 
    -101.706487745348, 
    -129.963507125787, 
    -174.564456409995, 
    -163.244905866941, 
    -163.64761607137, 
    -187.492392743956, 
    -141.182442108701, 
    -76.0154905105626, 
    6.03585458546053, 
    81.5708328943366, 
    101.75029199094, 
    65.8375477780152, 
    156.787766389325, 
    98.453572684414, 
    29.5361575733233, 
    -35.8689728087535, 
    97.1770893259263, 
    188.417690321955, 
    345.194143694702, 
    321.551790235289, 
    467.329255918901, 
    669.129455993582, 
    821.719159296078, 
    906.546971994967, 
    730.685497561606, 
    1440.11849285267, 
    1779.39034090972, 
    1407.19262977249, 
    827.701039996676, 
    453.83496789195, 
    1010.88724392232, 
    701.691578701629, 
    353.997875536163, 
    1026.26055058974, 
    283.932278491082, 
    65.3734192821475, 
    -3.60653161922729, 
    89.8235998410037, 
    -172.196971774771, 
    -324.511211151773, 
    -262.594957904878, 
    -189.124152904394, 
    -159.546982341223, 
    -180.717483761863,
  
    -2089.13472475263, 
    -1936.2034830433, 
    -1051.67128887796, 
    -440.176696743169, 
    -317.30097428308, 
    -215.353848073944, 
    -121.822686331002, 
    -161.844301608215, 
    -571.435845574765, 
    -973.231034786144, 
    -579.539147798851, 
    -196.443830972823, 
    -191.857694173046, 
    -33.1329517839743, 
    200.279083537094, 
    170.34467279684, 
    439.808106203495, 
    470.017514394352, 
    655.377013664631, 
    640.87448443918, 
    487.10400116804, 
    492.281871590609, 
    459.514772148175, 
    489.318888028819, 
    342.414272376698, 
    245.385772643137, 
    266.349812916652, 
    267.607078411277, 
    185.227120419766, 
    44.5464593702036, 
    -86.1365244567464, 
    -34.3859054470915, 
    -154.988350307555, 
    -210.995944991758, 
    -124.424284846358, 
    -156.383015125356, 
    -164.849531066912, 
    -187.163180162231, 
    -166.588333665991, 
    -76.4540409481134, 
    -2.71602086821249, 
    51.6216067845986, 
    91.9812117178265, 
    146.608560801353, 
    230.300571640289, 
    217.811405487316, 
    66.6128238366137, 
    83.0479976877262, 
    302.471010197451, 
    241.024193777616, 
    228.361489880125, 
    413.147360435393, 
    449.478605152912, 
    516.164805302294, 
    669.457330607621, 
    685.684919188566, 
    1237.05531498994, 
    1596.35687795812, 
    1585.61997052884, 
    1256.28287168633, 
    420.992488759618, 
    97.0578259386038, 
    912.392995973181, 
    1106.31142901413, 
    768.048707618156, 
    591.42113112976, 
    198.482157849251, 
    -105.107728774445, 
    -315.081520704247, 
    -199.718353591871, 
    -335.949654736151, 
    -274.9940633101, 
    -184.156485434742, 
    -130.376107266075, 
    -164.10775836291, 
    -193.744114659001,
  
    -1832.49055164845, 
    -1341.53857893479, 
    -594.783781677449, 
    -352.910879252605, 
    -298.506619290034, 
    -189.415336946357, 
    -139.997807241101, 
    -182.343354491077, 
    -534.161186423305, 
    -971.262760892826, 
    -367.640995734748, 
    -197.715141774826, 
    -149.392537998058, 
    36.5961106144067, 
    216.956579586425, 
    232.139692453894, 
    245.635089887082, 
    401.851508632887, 
    578.593335987872, 
    664.054225532898, 
    391.479268743636, 
    490.030511260166, 
    538.052939172556, 
    541.80226926387, 
    244.038836080843, 
    221.267309490003, 
    227.182349065116, 
    206.088055220856, 
    148.860300429324, 
    152.134261976031, 
    93.4966510231251, 
    -27.974536498744, 
    -67.4966155529561, 
    -138.858628696984, 
    -137.011180192065, 
    -172.460193354232, 
    -193.092489697498, 
    -195.99419268088, 
    -136.50048471218, 
    -19.5135720678562, 
    25.4627114480985, 
    92.550885273121, 
    143.770019883672, 
    155.104089531893, 
    184.575355867256, 
    230.424768065551, 
    104.81218078075, 
    -5.16527780573465, 
    159.37647290673, 
    229.754848499447, 
    268.284944876044, 
    448.267037732337, 
    450.401100338106, 
    569.952117005762, 
    813.001701679638, 
    1125.47798982046, 
    1776.39315611358, 
    1630.06594047247, 
    1514.70947050327, 
    1160.92295927964, 
    677.007161041107, 
    312.298186854325, 
    812.203698750972, 
    444.448963058491, 
    835.662284176133, 
    580.408890206232, 
    165.522750042852, 
    -261.114493138313, 
    -453.530756216701, 
    -408.028947917771, 
    -298.42713484812, 
    -165.288729190292, 
    -173.010301053858, 
    -192.170949290875, 
    -189.598461527039, 
    -195.553468638011,
  
    -1301.91036531079, 
    -626.19204658944, 
    -463.66018194047, 
    -289.445907567143, 
    -244.67512704437, 
    -185.856361032467, 
    -164.475407524579, 
    -213.961225973132, 
    -583.156317536799, 
    -734.231637345984, 
    -335.496537220304, 
    -117.609453579346, 
    18.7635006917289, 
    185.603466980135, 
    144.81739526046, 
    187.331240110409, 
    268.846617490421, 
    300.191502967313, 
    560.028026439843, 
    555.798443306199, 
    509.043459619947, 
    491.154126708744, 
    555.618252078202, 
    357.29204862195, 
    160.439128224286, 
    154.477483962978, 
    90.5002221826211, 
    84.2372983225515, 
    101.724135804683, 
    72.2516228648068, 
    48.6665155326924, 
    -24.1557619326057, 
    -82.9029122776572, 
    -205.858427711991, 
    -160.339141807257, 
    -211.528657904665, 
    -220.763275669777, 
    -240.238947066321, 
    -180.356252211072, 
    -35.83822882963, 
    44.3843768382528, 
    78.9994203726627, 
    119.031645645621, 
    132.405643616919, 
    160.686478814513, 
    178.6653899463, 
    104.924654098801, 
    134.133599707421, 
    -24.1018956020598, 
    81.2645982654738, 
    104.144568678779, 
    263.367544644089, 
    463.249074152042, 
    601.504519625981, 
    976.939922806931, 
    979.832581412222, 
    1433.83880126544, 
    1643.03022075794, 
    1367.18878537783, 
    981.387688503284, 
    398.792953980318, 
    106.850017102822, 
    931.449343340656, 
    657.23101879261, 
    606.059865069411, 
    160.408849609382, 
    -266.393779957548, 
    -188.276096727384, 
    -220.556587015262, 
    -242.557422924146, 
    -156.437794146052, 
    -167.822042676663, 
    -206.619320765855, 
    -209.097981498864, 
    -211.192663893321, 
    -213.362923809022,
  
    -740.44382375138, 
    -446.082098299818, 
    -440.231294638365, 
    -304.359841730132, 
    -209.965280282938, 
    -262.061082466187, 
    -337.140248455634, 
    -453.780144438367, 
    -431.390330507933, 
    -602.766683537908, 
    -184.986609282711, 
    -37.2251581966805, 
    -9.48293920486942, 
    156.82241207595, 
    223.16687287462, 
    360.494131385146, 
    290.313578205172, 
    352.526839957926, 
    269.559457894267, 
    276.433269804027, 
    392.693397436537, 
    182.155779867397, 
    282.758590668338, 
    204.152539476433, 
    144.288733234597, 
    106.397786732083, 
    78.942818891561, 
    46.4367538384863, 
    52.5567971797696, 
    -31.6171667083252, 
    -73.852339419914, 
    -59.8946221731816, 
    -107.285266865542, 
    -77.0685261740257, 
    -157.417106295219, 
    -214.912553539468, 
    -228.810032676876, 
    -218.696899085136, 
    -184.998390977353, 
    -98.2156543464702, 
    1.13259701686044, 
    -5.06800951422452, 
    63.5041805926255, 
    50.7419943521161, 
    159.699082305156, 
    205.023171759133, 
    194.400062016383, 
    157.771526458415, 
    56.9692374058033, 
    -2.33281299728877, 
    -165.174859257322, 
    175.355548296905, 
    223.673264459694, 
    344.610991508936, 
    388.400343793498, 
    604.90411749453, 
    808.365953597088, 
    1801.31675311833, 
    1515.50038126468, 
    963.419015591786, 
    447.238286618543, 
    14.3411756561783, 
    595.356435034602, 
    42.3392800894653, 
    122.63830418816, 
    22.8535851828745, 
    -262.913285113395, 
    0.47152666962746, 
    -171.536218048345, 
    -168.756507536061, 
    -86.6016548654409, 
    -151.751582951989, 
    -168.726587030682, 
    -177.417514341809, 
    -197.646478969066, 
    -196.213224539164,
  
    -608.301893740458, 
    -370.040270703904, 
    -416.97084066769, 
    -369.378418225057, 
    -481.464511209213, 
    -543.919680118029, 
    -679.214912252224, 
    -722.303171429094, 
    -467.805499163349, 
    -465.90319077512, 
    9.19381241008405, 
    36.5646785838084, 
    321.783084700651, 
    330.052217955553, 
    402.335665229721, 
    212.346162851553, 
    170.662447569486, 
    398.786045437563, 
    246.693289514351, 
    62.0023786196652, 
    190.02956110793, 
    181.685645170735, 
    69.7858358625594, 
    27.2707649708332, 
    89.0747867009676, 
    82.9529879378847, 
    24.3135003496257, 
    19.2610461958845, 
    -44.9821961179693, 
    -67.1478796475142, 
    0.924718004191147, 
    -43.0883896850133, 
    -196.900431007179, 
    -54.3547214767567, 
    -167.13510019061, 
    -198.755266178896, 
    -235.128236913734, 
    -203.646883634544, 
    -185.615529108421, 
    -153.951563372724, 
    -114.212971099947, 
    -60.6240037942653, 
    23.9342983397768, 
    76.4938123549217, 
    94.7743823183873, 
    174.743720318409, 
    162.910927596312, 
    185.069833106184, 
    66.5879118162859, 
    245.589740582303, 
    -109.310807252649, 
    -33.3407683064114, 
    291.530320674816, 
    341.83541575792, 
    461.233557415975, 
    974.951825644913, 
    1248.86389939328, 
    1269.27603689366, 
    1082.57618231522, 
    812.799334475866, 
    379.977617962219, 
    -82.6425007377398, 
    101.759522713443, 
    45.268106750584, 
    76.4093049720565, 
    -199.215078187283, 
    149.657411372412, 
    -82.9295898194016, 
    -200.963853419562, 
    -125.698250193878, 
    -127.565018018444, 
    -217.82908322376, 
    -238.817080573567, 
    -272.066369418736, 
    -271.948838420839, 
    -259.080238508885,
  
    -554.055136916618, 
    -395.574418250551, 
    -382.453151463661, 
    -439.704099512046, 
    -585.592489928174, 
    -725.23609855968, 
    -413.123341563561, 
    -407.329241172727, 
    -112.549838635313, 
    -89.1728549815224, 
    3.65528130745042, 
    125.836139957689, 
    303.194619041003, 
    280.075814088006, 
    309.721397113692, 
    289.730383011155, 
    214.077911221035, 
    161.54089736832, 
    219.13823927637, 
    182.067625052185, 
    211.838732910584, 
    174.568254092773, 
    84.8250425206321, 
    73.5180128370931, 
    144.567510070887, 
    98.0568250856901, 
    40.6387944888958, 
    5.08094635435545, 
    -45.2518026270768, 
    -69.5674645972825, 
    -77.6666361375206, 
    -205.300280888162, 
    -84.059391585601, 
    -73.5794165024967, 
    -119.46608536668, 
    -175.745444518855, 
    -205.669742917427, 
    -207.959472338003, 
    -197.057967671889, 
    -181.51768370198, 
    -132.202817748135, 
    -84.1631667050643, 
    -24.0049131107492, 
    63.8176693013894, 
    77.1797520513661, 
    150.984580696763, 
    249.639403310094, 
    321.061757351491, 
    227.65648914051, 
    56.3198968886248, 
    163.912853612611, 
    -99.0017238886079, 
    115.699915463018, 
    401.536644323676, 
    513.062087662411, 
    929.636099777993, 
    1278.52218255431, 
    1331.72843063372, 
    1086.37856103912, 
    911.12727162018, 
    -13.7191032551799, 
    -32.8274606967867, 
    282.079182394141, 
    -13.7064460727024, 
    -143.533550438663, 
    -82.5224498575724, 
    -3.17538475990403, 
    -128.464576540709, 
    -259.609449566013, 
    -260.19970467323, 
    -238.745970618153, 
    -305.792323480929, 
    -300.744087159433, 
    -326.635227946657, 
    -332.734096779134, 
    -349.077511974305,
  
    -519.240026480407, 
    -406.701189171428, 
    -321.890025887482, 
    -151.662970989307, 
    -134.218948732291, 
    -422.753108056627, 
    149.208499286908, 
    16.8551425770842, 
    249.656901646837, 
    31.9818685612783, 
    619.627296131641, 
    639.910899693063, 
    257.573727418708, 
    271.783937580243, 
    311.624001745414, 
    429.435532803765, 
    447.014619440674, 
    307.374401865722, 
    173.610123477351, 
    270.376775662549, 
    315.840067112699, 
    187.992921164962, 
    110.783891556111, 
    112.154470973427, 
    153.049813756483, 
    112.668934654415, 
    -23.02390700572, 
    -43.793360588933, 
    -93.775281236527, 
    -206.485807984833, 
    -134.664973549452, 
    -86.726472460543, 
    -53.2897037130198, 
    -101.078477618142, 
    -150.408404998523, 
    -165.718332034343, 
    -177.040595418795, 
    -181.379972009348, 
    -159.964410166724, 
    -157.400109657381, 
    -123.810326766327, 
    -104.664337687904, 
    -87.5348460484729, 
    -71.7572473278247, 
    93.5785338731762, 
    -16.8924843797772, 
    136.109402932084, 
    290.799342743893, 
    316.860982029862, 
    270.339592462692, 
    238.075160565863, 
    244.515305434735, 
    62.1120532837894, 
    150.186351436516, 
    263.01709764081, 
    524.732711334909, 
    752.289323761905, 
    1313.87833417355, 
    954.99081203892, 
    778.560009276064, 
    -177.265603581314, 
    96.9041399309702, 
    229.752430679824, 
    -2.03495989631521, 
    25.1915969128055, 
    72.9912156999989, 
    -148.043466020137, 
    -209.61175679787, 
    -293.800931612295, 
    -293.912522977036, 
    -275.325594586996, 
    -268.114663580097, 
    -249.304616223256, 
    -211.308884386786, 
    -208.033992818596, 
    -320.814675567128,
  
    -498.648953137713, 
    -422.177041232119, 
    -255.074587423616, 
    -56.666438268782, 
    127.943971494011, 
    60.9244753569575, 
    125.381830391662, 
    436.624580379031, 
    334.017291125636, 
    646.965690775127, 
    801.143717408051, 
    528.565873713137, 
    660.88926486606, 
    522.967557601674, 
    278.211205442969, 
    389.853772410086, 
    401.125810514239, 
    298.026690146691, 
    141.037067699539, 
    145.170374540305, 
    247.918482089495, 
    210.885439752064, 
    141.132863035128, 
    173.691891120236, 
    56.7318410793312, 
    24.5766568534978, 
    -30.2824108429749, 
    -48.9616620591348, 
    -130.71190093426, 
    -109.97614108061, 
    -136.238276965408, 
    -146.133237947676, 
    -134.020192076885, 
    -111.61134371592, 
    -162.487551645362, 
    -147.502443140592, 
    -151.4790336752, 
    -140.145071520918, 
    -145.73492234071, 
    -97.9792001185998, 
    -115.597410696485, 
    -107.035605613221, 
    -116.638963205951, 
    -130.420983666936, 
    -144.887580675081, 
    -139.274893662431, 
    1.51736934027445, 
    174.50118722307, 
    247.712809854233, 
    328.339571005553, 
    263.061541225181, 
    81.0527332755493, 
    281.31721614056, 
    341.214868487862, 
    103.989898631447, 
    240.250367043934, 
    270.020703254861, 
    549.828723864762, 
    808.369856198978, 
    188.732026936352, 
    -278.006697262791, 
    282.448648358785, 
    451.589156681578, 
    130.159209611297, 
    284.449834639924, 
    257.32597521091, 
    -136.016926552387, 
    -281.295734362798, 
    -236.555333431195, 
    -204.560964614253, 
    -223.219984817078, 
    -227.913379344534, 
    -220.298966302049, 
    -200.217806018347, 
    -187.764905088025, 
    -203.748191483211,
  
    -532.337211617431, 
    -400.910450259355, 
    -88.2260767398977, 
    474.53906682304, 
    181.6445625899, 
    390.828130707098, 
    509.478989869189, 
    670.39841781565, 
    829.682880269188, 
    817.615963550323, 
    753.345747935943, 
    531.549675423515, 
    562.234552765747, 
    567.22474168049, 
    471.885036647922, 
    398.655765131903, 
    315.896501654339, 
    239.113266392758, 
    157.011066387642, 
    140.049961786387, 
    183.227075818139, 
    204.427531194313, 
    149.629236061122, 
    70.9214065269806, 
    31.2807718994629, 
    -3.6288542599325, 
    -68.5601071360932, 
    -86.3307592940896, 
    -150.588484581481, 
    -132.073619690881, 
    -148.58557320709, 
    -178.328173185649, 
    -168.288985746839, 
    -271.758214431542, 
    -213.78686934596, 
    -177.175385138756, 
    -244.822839478495, 
    -201.595803031195, 
    -264.477348637341, 
    -128.256444187741, 
    -131.465927064218, 
    -80.3201228501675, 
    -109.437304682588, 
    -129.707432997854, 
    -182.067425978812, 
    -244.604436878662, 
    -116.228485186451, 
    23.5053870576476, 
    258.142771431473, 
    320.312610997865, 
    262.776635438037, 
    162.697883225771, 
    328.373198749506, 
    232.866275595122, 
    66.3636552011386, 
    371.220537439845, 
    99.554958259137, 
    439.542736301223, 
    316.350908233489, 
    -238.963957682971, 
    -227.170627831071, 
    372.08256573907, 
    495.180794146675, 
    352.932820297699, 
    357.478294364014, 
    296.515502233381, 
    -140.925452901962, 
    -191.393746716712, 
    -162.047783455415, 
    -206.519027801805, 
    -223.794497249642, 
    -234.734265503665, 
    -222.091177313485, 
    -208.641375393243, 
    -205.796352484727, 
    -273.670413125136,
  
    -598.637966279888, 
    -308.295871879859, 
    -19.907305399754, 
    488.765299114639, 
    506.149575783448, 
    497.883805589994, 
    250.649482336178, 
    805.770131434735, 
    882.621212112409, 
    634.533710073917, 
    748.28894536786, 
    653.700971007481, 
    560.780455158914, 
    554.605696281954, 
    530.151930062527, 
    383.326389727106, 
    249.518647701181, 
    201.801680414299, 
    89.8280694060192, 
    116.280548223858, 
    201.445205257027, 
    186.668990524992, 
    127.129308438915, 
    47.2348932846128, 
    -8.54387490219425, 
    -22.3156686648808, 
    -73.2476967868186, 
    -94.4081291121837, 
    -138.044437083792, 
    -179.118454857342, 
    -111.669310226953, 
    -81.7906326024828, 
    -147.037840350879, 
    -154.678441651056, 
    -112.575918527626, 
    -80.4264407387515, 
    -108.510455637736, 
    -131.677608277471, 
    -237.26037797789, 
    -196.183658595582, 
    -92.4307105618643, 
    -13.7524877460914, 
    -127.251133613328, 
    -113.201647096357, 
    -127.072995837298, 
    -138.776192234718, 
    -244.146276138666, 
    -163.655060342018, 
    152.697644717482, 
    286.153303639752, 
    310.150873908271, 
    244.845754476033, 
    248.487921602651, 
    279.942525019971, 
    274.39818125956, 
    612.315448534577, 
    173.061227616911, 
    293.1160212834, 
    257.571089506425, 
    270.484436289336, 
    6.43213883706811, 
    271.212886250706, 
    228.033455228212, 
    97.0205156127573, 
    65.5593350452892, 
    -0.477041602942018, 
    -189.989742603708, 
    -173.898059785165, 
    -198.72421198436, 
    -204.681709407024, 
    -245.864216673147, 
    -214.676467088141, 
    -201.622336435692, 
    -263.710352430954, 
    -304.497114102491, 
    -309.351789532156,
  
    -636.051773413031, 
    -210.619206824735, 
    209.840964660131, 
    306.22815211809, 
    320.537015000752, 
    378.165139705587, 
    743.870285820193, 
    813.368462967306, 
    632.718064055061, 
    666.586784362791, 
    599.977466365392, 
    584.66918542911, 
    595.272940094233, 
    539.415441002584, 
    561.085144974216, 
    365.443945638008, 
    186.100702119166, 
    100.414381749152, 
    138.447469888585, 
    200.871471005619, 
    207.08832050678, 
    178.424345121138, 
    132.620016163167, 
    60.0637341805829, 
    -22.5258720336277, 
    -43.0211121259054, 
    -80.1781104601511, 
    -137.854415953359, 
    -174.353856391095, 
    -176.698881219776, 
    -141.117053045805, 
    -130.552571648046, 
    -170.119128901106, 
    -109.542946024143, 
    -60.7658746506832, 
    -104.54052792044, 
    -122.202308660124, 
    -147.037704537189, 
    -193.196321083742, 
    -153.516066009758, 
    -51.9483249713425, 
    -23.2977095798309, 
    -20.530512795337, 
    -122.461532239286, 
    -74.5170296565413, 
    -61.6979924908935, 
    -131.185892115781, 
    -100.375206358888, 
    96.6160061292664, 
    264.974797205053, 
    311.504193428782, 
    246.877269114787, 
    353.838544360734, 
    128.558513926358, 
    320.328741327779, 
    299.631020779837, 
    147.741620182331, 
    619.287706595124, 
    751.700256586877, 
    574.095772908755, 
    180.481487094752, 
    370.333994097567, 
    59.7598657997838, 
    40.0516383154099, 
    -111.178456928001, 
    -142.618885505908, 
    -188.518436634793, 
    -179.07928322838, 
    -239.480687563257, 
    -208.329420320398, 
    -206.204281126667, 
    -217.902492743191, 
    -226.008085368329, 
    -280.139070307955, 
    -295.121257235195, 
    -316.5056959966,
  
    -579.168850273992, 
    -114.296344923681, 
    11.244330762757, 
    -107.667592851202, 
    128.677958468179, 
    345.498992894298, 
    671.608576553541, 
    679.184820168763, 
    612.633118419067, 
    483.054990646686, 
    566.913237987144, 
    604.867284623132, 
    577.879555995893, 
    517.150571671472, 
    570.80827723692, 
    357.575723735642, 
    163.527662390424, 
    154.621816818822, 
    307.812336899265, 
    299.315221976592, 
    204.429717684379, 
    114.541326600787, 
    79.3217504529107, 
    53.3340829932533, 
    -32.1345480123802, 
    -63.5095553382116, 
    -80.581042809823, 
    -65.7325519239248, 
    -147.954173879419, 
    -180.610615705723, 
    -188.223551670088, 
    -112.534864730023, 
    -104.31254898554, 
    -74.0783377355853, 
    -42.8540959037839, 
    -92.7320327769473, 
    -102.757962793946, 
    -51.4572989628262, 
    -16.9100148375461, 
    19.9152433548183, 
    -32.2730211688323, 
    -48.1435511947884, 
    -29.8851850969931, 
    -122.085144453058, 
    -26.917730176434, 
    7.69940017752885, 
    -6.12474238425226, 
    -38.3044840731511, 
    29.5886639056247, 
    120.717357183756, 
    260.145785499393, 
    179.806140750147, 
    173.918404821584, 
    -48.0166454130976, 
    -69.0316983155737, 
    90.2199628131501, 
    442.78804440728, 
    652.288275373744, 
    682.834379241018, 
    464.089981698506, 
    135.091295448151, 
    337.87395033884, 
    386.407358923515, 
    210.711872171301, 
    -50.7691869383284, 
    -130.09121751278, 
    -120.787389410305, 
    -249.47294664757, 
    -282.387948710068, 
    -318.703245588005, 
    -277.710145303143, 
    -264.542785537737, 
    -276.025833625409, 
    -300.063414865219, 
    -343.532617686445, 
    -329.558557550958,
  
    -492.354380198582, 
    -274.646384129206, 
    -110.70995246443, 
    297.75850220838, 
    716.102515157634, 
    683.129422793335, 
    723.198257779479, 
    508.384885918242, 
    382.788497766747, 
    450.549068045114, 
    444.304539957077, 
    577.019780183558, 
    543.980657622369, 
    561.291620226751, 
    549.560506728836, 
    325.028097312901, 
    242.459705673168, 
    422.101428613952, 
    342.024120065961, 
    205.045139430219, 
    154.487970782553, 
    96.6717345706545, 
    79.1007334740133, 
    14.0316956320905, 
    -90.63538104289, 
    -64.6079070698903, 
    -74.8574464569427, 
    -64.9316017550292, 
    -99.261299011555, 
    -151.640040310072, 
    -234.309046945007, 
    -133.975944953696, 
    -118.997680500668, 
    -100.799659935118, 
    -73.4155174321586, 
    -115.117810349715, 
    -119.602552749274, 
    -31.0377684432474, 
    -116.298966325546, 
    -88.9043736441822, 
    -104.570280297207, 
    -68.7676408058576, 
    -30.2191372465036, 
    7.66725057290236, 
    34.9669732414741, 
    62.5821909562737, 
    31.7361581517754, 
    -27.0244755643487, 
    33.8933118454968, 
    -41.7395410780695, 
    239.459247452414, 
    290.180072100939, 
    256.070223884111, 
    58.2573158460705, 
    -155.499320255548, 
    -175.111748271401, 
    228.880795238539, 
    849.886870175962, 
    421.132725735922, 
    377.029989317308, 
    136.602861669994, 
    25.4102612978107, 
    48.0721625012189, 
    -21.2580306238327, 
    -36.2506209754725, 
    -52.7249240146418, 
    -223.934171595474, 
    -328.159078783846, 
    -316.313846037076, 
    -286.793664772059, 
    -265.259120441364, 
    -265.41341927711, 
    -260.1078744805, 
    -384.897075025127, 
    -439.356409570541, 
    -391.240131737004,
  
    -433.699130319934, 
    -610.344434919713, 
    101.636076960027, 
    222.588309466386, 
    595.252131599868, 
    669.2589145844, 
    257.272659188556, 
    624.788901052441, 
    498.513999622842, 
    613.002205381989, 
    174.335810446658, 
    508.454532008155, 
    566.513206481933, 
    591.639863615474, 
    497.840901634328, 
    284.113359500421, 
    383.276525307346, 
    442.959599839878, 
    303.995257062578, 
    196.514753439924, 
    135.281456283065, 
    70.7950398022223, 
    25.2524242708146, 
    2.97966366567418, 
    -56.6426498481424, 
    -39.0437097597495, 
    -48.223957963113, 
    -55.5107318620802, 
    -92.6638707911718, 
    -89.0331977713943, 
    -115.23855084294, 
    -103.774041253801, 
    -145.536204674477, 
    -135.92840455174, 
    -87.4646170296837, 
    -118.614299133404, 
    -150.825823071556, 
    -8.37586295885029, 
    -30.5785646753624, 
    -26.3610780694305, 
    -56.3859750746603, 
    26.2757031154335, 
    42.0494700396584, 
    49.42573133962, 
    59.6744299719873, 
    44.8792130784245, 
    12.7075506163074, 
    -40.6502865831887, 
    71.6153271390518, 
    172.019019657656, 
    73.4012769798411, 
    178.459365481621, 
    135.260614896006, 
    -59.1321233416163, 
    -244.455946143772, 
    -293.130991488261, 
    47.5728403331199, 
    561.906416274667, 
    192.289978620325, 
    55.0508823202525, 
    11.7803740787055, 
    0.382459166800635, 
    36.629368613306, 
    -63.5932704774649, 
    -136.293236827532, 
    -250.835129723976, 
    -362.948388769272, 
    -386.688934052778, 
    -354.987439577417, 
    -340.143679628448, 
    -305.56137234046, 
    -279.552974863256, 
    -246.96777943294, 
    -353.50067756371, 
    -448.347870565072, 
    -370.453616784106,
  
    -333.032085113269, 
    -859.072049259475, 
    180.760944172095, 
    654.064731943907, 
    702.533688535598, 
    133.118773081251, 
    420.521079357058, 
    -425.631331039038, 
    -111.926681315677, 
    313.683169385215, 
    212.661626527461, 
    594.397324736152, 
    679.587234616679, 
    630.385998306189, 
    521.713248394904, 
    406.936329460359, 
    441.621289499931, 
    340.536284554577, 
    109.906049085489, 
    92.4709489956936, 
    130.626202492538, 
    73.706399325961, 
    11.0761441539679, 
    -55.1954089716861, 
    -13.382785678043, 
    -39.6839442672284, 
    -103.61667182598, 
    -71.9759418652022, 
    -87.6347158716078, 
    -46.0487552030886, 
    -5.61456169513346, 
    -50.0978809850075, 
    -135.854877259403, 
    -143.093045591373, 
    -85.6812129175547, 
    -113.35578400504, 
    -97.1911958713676, 
    -40.6794702395352, 
    -33.1337148398342, 
    -9.38213145165695, 
    -45.3153548021741, 
    18.9960105642591, 
    36.7174051093623, 
    21.2651607860768, 
    31.3214455395768, 
    39.3109113729546, 
    40.9231612252501, 
    91.2592257235935, 
    211.943700625943, 
    111.689757567104, 
    85.0657308883932, 
    173.538104577404, 
    115.208690354962, 
    239.534716658472, 
    -173.472288911316, 
    -322.199924678311, 
    -47.0958619155053, 
    743.320245561248, 
    570.64409420445, 
    -75.3521650050985, 
    -19.1906611914064, 
    -18.5356339260267, 
    191.341061136081, 
    -119.377209178546, 
    -253.882326589588, 
    -410.83130202769, 
    -436.800232258249, 
    -401.831229377569, 
    -414.931148358181, 
    -376.358552127509, 
    -346.431405314138, 
    -231.109427839748, 
    -243.815180689864, 
    -330.983669456148, 
    -284.543899924863, 
    -293.599087953298,
  
    -262.792762685865, 
    -836.24685471588, 
    -636.944602124786, 
    -319.283553583791, 
    -706.409588513666, 
    -527.046228497961, 
    54.4334514367042, 
    619.449954999396, 
    407.365330306327, 
    528.848726637824, 
    576.781746534327, 
    635.252290279308, 
    608.671830428275, 
    620.606394768828, 
    569.517896910665, 
    483.3637323497, 
    425.608454496035, 
    296.948829492822, 
    120.065206274609, 
    161.671559497198, 
    136.877486255642, 
    55.5575862491513, 
    34.2443507267674, 
    -10.5318668428608, 
    -4.91249297133755, 
    -62.2722949901614, 
    -172.298829233525, 
    -109.387400698689, 
    -90.5733227628337, 
    -20.4967287590629, 
    -17.42885058551, 
    -27.9720609938307, 
    -116.402266933826, 
    -111.227114336753, 
    -103.5732877129, 
    -89.2988843330468, 
    -76.6640049420698, 
    -62.9838735333746, 
    -47.9883893804345, 
    -104.472998697038, 
    -96.4026795907343, 
    5.77229041208179, 
    16.7201015325829, 
    -21.9199788938844, 
    11.17936393068, 
    50.0246623424784, 
    63.0807109888314, 
    168.797594963237, 
    213.460532813162, 
    154.23800652772, 
    95.5902177911049, 
    156.415593150481, 
    16.5960385704631, 
    -21.1919066709793, 
    -283.32710356675, 
    -396.030883507123, 
    -104.218312625655, 
    477.384232148332, 
    551.431951251559, 
    301.86510325279, 
    -24.1682202175247, 
    -26.1122327582436, 
    1.30421413359271, 
    -140.428609574629, 
    -255.60218875112, 
    -411.154145389227, 
    -338.571853150708, 
    -270.353212081034, 
    -306.719057350114, 
    -324.995160170123, 
    -294.841890162074, 
    -180.850321762241, 
    -225.765259619924, 
    -251.041070034629, 
    -260.048829835846, 
    -159.288802434189,
  
    -403.308528652384, 
    -332.086484851386, 
    -248.344904961501, 
    -1.90214010007788, 
    -23.206784167995, 
    348.8682748895, 
    438.573988757488, 
    548.108517850765, 
    933.847776398011, 
    718.810390066596, 
    747.201061321401, 
    680.084691627561, 
    650.50785907946, 
    601.478451676491, 
    539.829116060911, 
    496.768278359031, 
    415.972366986588, 
    283.38346872618, 
    155.441204013377, 
    177.106572596516, 
    129.607413082613, 
    13.2252685656933, 
    6.90258511894485, 
    38.7420040239552, 
    -68.303724626944, 
    -138.917564484999, 
    -93.6018960809655, 
    -97.1958841748892, 
    -46.0963426752274, 
    -8.23629330413902, 
    0.669579626064979, 
    -2.33479775813898, 
    -92.4968999881883, 
    -38.2846384280735, 
    -46.5241338363006, 
    -40.1327361574632, 
    -48.9551187981954, 
    -27.6992806726175, 
    -39.0633104053086, 
    26.8694704525409, 
    -32.9836336741393, 
    -17.3879303108536, 
    -17.6383949970753, 
    9.83265131565211, 
    32.1736560556689, 
    72.5180135878578, 
    179.679984093782, 
    216.388494410416, 
    224.622617796314, 
    150.360612459172, 
    99.0474668750583, 
    64.0516314874971, 
    15.9960944130091, 
    -143.4567914196, 
    -207.647423670513, 
    -316.914536970594, 
    -275.705427095042, 
    -34.5499214234366, 
    -69.7002759871661, 
    -19.105590385736, 
    -12.670694661365, 
    12.3990206818282, 
    83.9296156827375, 
    -151.800696573761, 
    -303.385714668711, 
    -243.469621173472, 
    -114.530195053585, 
    -194.700497566386, 
    -226.96518182701, 
    -238.383070156528, 
    -201.693861740299, 
    -218.428630256439, 
    -228.515183202096, 
    -258.333025339603, 
    -245.417540512853, 
    -229.976870245257,
  
    -474.947794654735, 
    -293.229476014548, 
    32.0613178411119, 
    -91.682439463403, 
    -57.9335988451628, 
    472.018090742551, 
    505.654974404529, 
    708.357361463523, 
    738.509243186616, 
    724.194139521169, 
    705.050091742398, 
    624.737244575048, 
    524.569037041232, 
    576.801881147258, 
    512.934357031194, 
    425.057591057036, 
    351.476393499939, 
    238.86306805413, 
    136.578317142411, 
    80.4772806915128, 
    107.489482627604, 
    80.3666470357844, 
    -15.0414486714999, 
    39.671123124451, 
    -22.8956127884922, 
    -33.5358862011847, 
    -61.0722337927811, 
    -43.8509128219183, 
    19.3033984519078, 
    74.6021763885969, 
    -49.8195728067624, 
    -2.81372219016905, 
    8.41533548441205, 
    15.9021654218491, 
    38.3606030671368, 
    -15.1723043898563, 
    -50.4007668196139, 
    -33.239046962905, 
    -52.2404160189865, 
    -6.4448943138771, 
    -8.23628621045099, 
    -1.07693246058686, 
    -37.9875721952804, 
    42.2755225022451, 
    48.6397303792694, 
    55.1470357162295, 
    169.409341780094, 
    225.308241661559, 
    218.094103487448, 
    149.447859816428, 
    155.438321793867, 
    148.790144761222, 
    -31.8326137786761, 
    -204.665905707894, 
    -168.584997497506, 
    -243.923459342451, 
    -225.292551429382, 
    -291.56930896977, 
    -401.965292098672, 
    -494.725590064015, 
    -107.450812089351, 
    1.32668929183918, 
    28.3239738524658, 
    -250.781971375061, 
    -305.399077647209, 
    -128.501614854687, 
    -68.0606210586875, 
    -122.654573432007, 
    -173.923478439435, 
    -187.241052328538, 
    -184.782519484687, 
    -182.718882927035, 
    -196.383856050378, 
    -225.996477306489, 
    -218.805975759149, 
    -273.14939344263,
  
    -507.481038032701, 
    -204.904978996697, 
    -153.129179062796, 
    -106.476538335623, 
    89.1678126995581, 
    573.547607823419, 
    548.316658669328, 
    641.364604740633, 
    679.50484360613, 
    684.633560180668, 
    606.452187942902, 
    598.55132117704, 
    483.977858843486, 
    538.070531642182, 
    474.100867242587, 
    357.991011389959, 
    287.245053401318, 
    207.842709956751, 
    107.806033941827, 
    72.8880681532364, 
    117.153121746398, 
    46.1571669167381, 
    31.4952609456269, 
    39.0031643538566, 
    43.0086107617126, 
    13.219144797139, 
    0.126860343329099, 
    38.7527491899526, 
    57.6782860857378, 
    151.512568547504, 
    -151.784480710045, 
    66.3810915546525, 
    112.715913593169, 
    116.855214332547, 
    131.081905448291, 
    142.577433172829, 
    38.521537035872, 
    -34.7316703331832, 
    -39.0228658341878, 
    30.5273985694863, 
    55.6867630553792, 
    -7.48395682449168, 
    31.5336754682506, 
    22.5215703853036, 
    62.0899158810988, 
    93.6430321295092, 
    147.572791410321, 
    226.212177479522, 
    227.296374426711, 
    188.100377788737, 
    139.273588825581, 
    38.1124983277735, 
    -56.3971762966868, 
    -132.589739443872, 
    -81.9687297501692, 
    -87.1464202788442, 
    -195.311062087669, 
    -190.885649351108, 
    260.235771422712, 
    433.714921363933, 
    21.9135480917638, 
    -41.5116021310107, 
    -31.8612500709479, 
    -289.200953230478, 
    -261.105458713456, 
    -70.9992581065261, 
    -97.8586327978905, 
    -97.4784760640696, 
    -198.927421668074, 
    -191.519259579905, 
    -184.423655846352, 
    -200.092166597339, 
    -196.112196462018, 
    -212.37596214098, 
    -197.845245542878, 
    -270.663524689625,
  
    -661.97929941927, 
    -297.004764172425, 
    -191.433173586513, 
    -79.6270280466368, 
    306.967501402167, 
    738.25992140818, 
    860.077850239274, 
    642.092967717938, 
    661.218201982214, 
    753.693993913367, 
    640.229079909714, 
    360.616034927454, 
    446.071129891801, 
    481.690517015447, 
    396.871748203393, 
    321.614402736822, 
    233.732721044662, 
    164.999098129529, 
    93.8475773043488, 
    86.0201013229731, 
    14.738866601452, 
    48.1911758196446, 
    39.2123147829918, 
    60.7721008944752, 
    61.317197829585, 
    65.4187423667607, 
    48.7458432625816, 
    79.0244509962878, 
    131.249910719851, 
    195.311413686994, 
    -137.381225674577, 
    239.247521570255, 
    139.847537348278, 
    120.204004326166, 
    182.590277121823, 
    212.755936181559, 
    103.073676406202, 
    -1.71057497270319, 
    8.84797072116894, 
    63.1663906181779, 
    132.567095364595, 
    117.191633967776, 
    95.6026160965306, 
    115.955153087219, 
    151.403596147578, 
    178.29836084808, 
    203.30148788529, 
    266.51937371112, 
    307.987209610549, 
    309.084639084699, 
    275.615122078514, 
    163.146075491141, 
    55.520819724339, 
    -37.7764350972812, 
    64.8440847396855, 
    120.824928856111, 
    -73.4676354393375, 
    -426.051801722101, 
    785.320873341663, 
    504.148766909576, 
    139.780159064392, 
    -108.644850991474, 
    3.63970588009128, 
    -218.544265535618, 
    -68.9705113670456, 
    -62.465100846926, 
    -55.0237362029704, 
    -160.72016912078, 
    -190.589599427824, 
    -186.738291346346, 
    -194.671060406214, 
    -227.459638065881, 
    -220.144744433054, 
    -250.039318804511, 
    -244.809190871869, 
    -295.137966946285,
  
    -650.238868653574, 
    -601.332633707318, 
    -345.630265969578, 
    -149.460056185321, 
    474.39784340255, 
    942.968809574208, 
    717.12232196291, 
    509.929595421837, 
    546.377434990041, 
    480.033589708044, 
    565.1902629942, 
    445.075272106244, 
    160.641115391508, 
    411.75135765631, 
    249.850186419514, 
    221.875657388104, 
    150.790465745787, 
    86.9063711748411, 
    61.521068692608, 
    40.0798391895358, 
    51.9419725531293, 
    66.2597920427394, 
    78.4880800033603, 
    55.0284577216975, 
    49.3921490724784, 
    107.210561914647, 
    98.9038991949459, 
    133.98188231747, 
    210.529599088304, 
    314.168794693899, 
    -24.4029852325434, 
    151.601799956361, 
    124.206435164038, 
    105.557037228566, 
    210.272739361275, 
    139.599509677054, 
    125.982843407591, 
    52.2234857026296, 
    1.51810689706008, 
    86.6371949004703, 
    266.572986402011, 
    281.063485785267, 
    147.987968299583, 
    185.151361574385, 
    166.243390065158, 
    190.143856659449, 
    270.500275602266, 
    324.606422018498, 
    361.021372433072, 
    404.6770415226, 
    436.220098305389, 
    354.935952766478, 
    320.954881324211, 
    59.8118258772075, 
    81.6862611952184, 
    201.589418972995, 
    141.972857959056, 
    -24.8846108466738, 
    -155.248038201155, 
    16.0495427551894, 
    -48.2463183990394, 
    -135.4025218938, 
    -197.930247335658, 
    -128.588134344854, 
    -49.0090826425413, 
    -50.0532548761315, 
    -78.3475807879833, 
    -112.266492760328, 
    -267.867876700033, 
    -282.794899772824, 
    -250.753165822813, 
    -212.622148345059, 
    -257.664174992987, 
    -204.19379164684, 
    -238.112044209463, 
    -307.360380132147,
  
    -596.712761728387, 
    -665.375577424702, 
    -677.183570861816, 
    -403.638182790655, 
    -42.2585956673877, 
    438.268328616494, 
    431.557578438207, 
    353.296443336889, 
    337.472434997559, 
    315.236446380615, 
    340.846323113692, 
    263.321685188695, 
    284.984640924554, 
    238.049924850464, 
    83.4608924765336, 
    58.3466552684182, 
    63.6377880196828, 
    -12.7775589729609, 
    0.626644556263556, 
    49.0243964697185, 
    68.5737583009822, 
    208.549541573776, 
    76.7998156798506, 
    36.5747619930066, 
    -16.9242688056672, 
    40.2908269480657, 
    140.566414983649, 
    189.570339002108, 
    252.178823471069, 
    272.433590537623, 
    -29.1812480625331, 
    187.717585312692, 
    143.666061501754, 
    87.3123190528467, 
    130.977451625623, 
    146.788390912509, 
    225.654082850406, 
    109.053473924335, 
    93.3320743661178, 
    52.9940614951283, 
    209.885619715642, 
    325.077346400211, 
    192.862276579204, 
    92.3126645339162, 
    148.611090609902, 
    238.040080923784, 
    304.831702382941, 
    364.181953430176, 
    405.965842397589, 
    449.491364127711, 
    485.902560786197, 
    468.654064981561, 
    441.720090364153, 
    5.76858553133477, 
    183.725795545079, 
    439.815229917829, 
    508.163236316878, 
    634.277794285824, 
    102.64456991459, 
    13.319924122408, 
    -107.022936820984, 
    -181.102675186961, 
    -201.628659599706, 
    -121.484992529216, 
    -44.5057888532937, 
    -54.6753153299034, 
    -101.331889152527, 
    -112.686148342333, 
    -230.452665328979, 
    -190.567063080638, 
    -363.475929461028, 
    -307.372620632774, 
    -212.179993880422, 
    -190.440703040675, 
    -264.862432178699, 
    -332.736596559223,
  
    -206.560856907792, 
    -328.89430820341, 
    -632.349982241367, 
    -598.887376210724, 
    -401.860506307639, 
    -83.087481089829, 
    -63.1387031038306, 
    -94.8510451710976, 
    -76.4597446381854, 
    -125.397805254511, 
    306.870134953822, 
    61.0422151198174, 
    8.58025908490144, 
    -121.20231167066, 
    -79.7055020604663, 
    -98.8263465955037, 
    -106.748483790262, 
    -71.9704801350131, 
    -56.6814170166734, 
    21.1560139513232, 
    290.464557154315, 
    290.567179894527, 
    62.7631716140829, 
    -12.5289878251839, 
    -70.0087251727287, 
    -131.39595916904, 
    2.62584239251133, 
    131.889913048484, 
    180.362345107058, 
    -4.86754315644467, 
    226.240965681942, 
    248.858777019505, 
    178.502690382528, 
    245.455138058038, 
    296.042222504652, 
    198.135281713385, 
    221.708992918555, 
    266.551288824733, 
    333.704866973177, 
    138.083218970731, 
    156.695011552212, 
    423.285305864733, 
    215.963365345492, 
    167.498848580834, 
    168.259283486566, 
    269.902318672531, 
    360.290169723357, 
    423.659245673647, 
    451.315554483207, 
    589.901677224565, 
    475.039754976484, 
    459.424314612103, 
    323.047575866252, 
    192.781880094118, 
    406.346911153763, 
    303.083685453106, 
    674.402745852417, 
    688.888600399619, 
    43.2108697116975, 
    566.474359811349, 
    480.037923452964, 
    -196.690905238853, 
    -202.605672274565, 
    -120.526247001041, 
    -51.2370668440088, 
    -128.350057837946, 
    -140.980622271274, 
    -147.806729534572, 
    -278.031060446284, 
    -270.505404768171, 
    -232.199431471701, 
    -199.755402143164, 
    -205.176028062622, 
    -214.188090859442, 
    -286.886781032516, 
    -361.01464375136,
  -200, 
    -200.006284292975, 
    -203.943994874516, 
    -448.001920198139, 
    -403.286216351379, 
    -394.286617830112, 
    -416.521434143169, 
    -343.45507125171, 
    -311.888671892087, 
    -282.535514750379, 
    -256.331185925048, 
    -311.685360245315, 
    -325.722665336071, 
    -376.302739116674, 
    -271.853566762448, 
    -102.07830654627, 
    -205.720237078352, 
    -218.217744607274, 
    -138.660071333472, 
    323.083550310084, 
    561.507260987901, 
    324.539096968972, 
    170.633251587461, 
    -65.3819642077638, 
    -171.176014125948, 
    -120.440473731661, 
    89.8819090874174, 
    334.965615608925, 
    117.346840441862, 
    325.416985463723, 
    384.57701745626, 
    191.516375119849, 
    220.303297036442, 
    487.770446375797, 
    443.612584283877, 
    287.901195462047, 
    354.662062569135, 
    359.140535083356, 
    390.465079488039, 
    226.560548139446, 
    254.393071613548, 
    284.71047392671, 
    137.766272614276, 
    102.198761500009, 
    168.135185980717, 
    286.700401325377, 
    444.651981802297, 
    530.132872723519, 
    498.467288633477, 
    602.24879963908, 
    708.195210515585, 
    302.601787447527, 
    368.465792212747, 
    130.207226629354, 
    345.889380041723, 
    462.111049882777, 
    206.742238464441, 
    695.172233590088, 
    64.9428766524002, 
    553.094056487213, 
    520.617359421946, 
    -169.902480818524, 
    -201.899013055799, 
    -98.5795121561367, 
    -69.2236042716874, 
    -170.70915981797, 
    -167.720226653079, 
    -253.230473132844, 
    -201.007505739389, 
    -194.348613706975, 
    -169.076341524369, 
    -197.450894226553, 
    -209.857842232853, 
    -303.403412091639, 
    -355.086713049741, 
    -703.410645855502,
  -200, 
    -200, 
    -200.703916133184, 
    -200.197205160126, 
    -202.047797120832, 
    -395.904212259632, 
    -306.980169294129, 
    -225.362671947159, 
    -187.924909657887, 
    -194.429100523603, 
    -209.536091675283, 
    -196.519199672498, 
    -193.789331476739, 
    -206.149819044089, 
    -215.549162852937, 
    -180.311603580316, 
    -202.420558673137, 
    -110.926075645948, 
    441.765372785716, 
    414.655552004378, 
    462.801704423825, 
    501.022742088806, 
    -56.8790556964351, 
    -176.249940167349, 
    9.38142229808705, 
    166.815871121503, 
    227.523639288086, 
    286.314378693548, 
    261.949171796758, 
    408.564225657123, 
    512.519249551908, 
    482.435473122762, 
    350.077350097436, 
    440.823639270573, 
    366.173949016302, 
    462.854522265085, 
    466.432687996484, 
    530.809363340611, 
    453.425577396508, 
    302.94690467262, 
    443.355975852704, 
    336.821863928408, 
    259.945431938899, 
    181.00477927743, 
    167.255007533451, 
    349.353773918026, 
    508.167384088908, 
    627.041620619754, 
    718.20205482577, 
    790.700719553573, 
    720.146995006189, 
    543.602473097713, 
    432.746160680209, 
    197.911114608318, 
    493.943708182717, 
    695.19187792258, 
    468.792146086821, 
    646.371360936868, 
    367.296933506267, 
    -46.6049028692434, 
    61.9872524436543, 
    -212.065644365678, 
    -207.516573915556, 
    -53.6816024539981, 
    -172.174741342381, 
    -192.535335970085, 
    -263.837706789058, 
    -236.861137116743, 
    -173.794840565988, 
    -176.845867142031, 
    -172.042383977841, 
    -196.749188742472, 
    -197.938770774765, 
    -412.776481568615, 
    -964.130864193572, 
    -1419.34386123709,
  -200, 
    -200, 
    -200, 
    -200, 
    -210.140894226638, 
    -328.203335506784, 
    -220.280254129065, 
    -217.947709229865, 
    -200.59402180252, 
    -196.038586839717, 
    -194.198567092485, 
    -166.650299082945, 
    -114.740938572173, 
    -103.289606114651, 
    -105.557237186197, 
    -129.960009276933, 
    -5.17252917786105, 
    485.931147080921, 
    411.738226519987, 
    444.052076764763, 
    451.879760191128, 
    227.219864575083, 
    -356.38219477108, 
    -211.927902328471, 
    305.119321415166, 
    508.85809016468, 
    469.548547242819, 
    324.415952834145, 
    238.708445406975, 
    515.125558171802, 
    530.285598797601, 
    308.455863694194, 
    439.766694999088, 
    399.568093627725, 
    545.951449685775, 
    506.796730857413, 
    463.019123649811, 
    641.568163462742, 
    591.898711534524, 
    511.908593121195, 
    580.120321643315, 
    487.465341390714, 
    577.21008492157, 
    532.30096911423, 
    323.875672313695, 
    169.212354019268, 
    373.479208041679, 
    608.522086285531, 
    694.73199879816, 
    794.171745377186, 
    872.687779092309, 
    612.124087808912, 
    441.044675829161, 
    399.497158528974, 
    371.460923890117, 
    780.388106402734, 
    565.241225615309, 
    491.523911291382, 
    815.255515932638, 
    324.870837682574, 
    508.89487122368, 
    -137.668196624768, 
    -205.181692202441, 
    -98.1670676067995, 
    -94.2364195260863, 
    -132.458521461701, 
    -202.871491817717, 
    -214.195150597499, 
    -205.922193369166, 
    -197.593083957275, 
    -201.922086252211, 
    -304.942339881138, 
    -434.094570873301, 
    -670.740009004573, 
    -1525.89787618845, 
    -2001.8980746894,
  -200, 
    -200, 
    -200, 
    -200, 
    -261.697509616112, 
    -200.162301303825, 
    -200, 
    -247.882089213321, 
    -230.881128813091, 
    -225.201845209649, 
    -202.007432568113, 
    -188.465781676409, 
    -132.500566684386, 
    -138.259390597115, 
    -90.8878683824956, 
    45.5535759046138, 
    255.61351070746, 
    244.429387708794, 
    392.404405860858, 
    342.812650229868, 
    310.696558769712, 
    -141.991794470848, 
    -153.980452750584, 
    373.757991876209, 
    501.051304910112, 
    473.402026241598, 
    451.205084323348, 
    502.743473394721, 
    269.331439403778, 
    617.176353941573, 
    478.72090255293, 
    238.8265727984, 
    136.238536616856, 
    553.55181075691, 
    627.022171251184, 
    463.087757448065, 
    453.626502845484, 
    613.437760484447, 
    681.571900840836, 
    635.49891223459, 
    629.364559630666, 
    703.293262930227, 
    606.876875028363, 
    605.161768581137, 
    530.35996590216, 
    210.875519268721, 
    203.697431888985, 
    410.117947679882, 
    643.419474243985, 
    747.0541590555, 
    693.693720100972, 
    682.258828209066, 
    656.361356177764, 
    648.517151075406, 
    187.509736164691, 
    905.107191335717, 
    618.615224114175, 
    553.147951085519, 
    205.848586322741, 
    6.28907493941707, 
    552.321754686235, 
    -45.4625028245017, 
    -232.785381712278, 
    -166.846074543234, 
    -151.387138215051, 
    -125.469593055571, 
    -123.536694344053, 
    -122.507885746031, 
    -204.437930528955, 
    -201.951853387967, 
    -280.594273021482, 
    -358.525284655016, 
    -591.359882119789, 
    -1357.22242926484, 
    -1831.25215866585, 
    -2160.74800924918,
  -200, 
    -200, 
    -200, 
    -200, 
    -200.457396333188, 
    -200, 
    -200, 
    -200.26142794875, 
    -218.550195758046, 
    -206.605610421363, 
    -202.892223821642, 
    -230.078549441672, 
    -212.288730226199, 
    -217.908387879375, 
    -103.486305708848, 
    324.038829517258, 
    467.855559751674, 
    555.169344928737, 
    648.147211277739, 
    219.373770422256, 
    417.097822631458, 
    -159.525525541616, 
    452.567991739433, 
    341.821369747828, 
    492.981864497749, 
    620.306412537715, 
    680.865325987541, 
    602.596239309961, 
    393.646396636964, 
    604.071754720416, 
    507.63841470118, 
    -245.271168763267, 
    361.176027693114, 
    500.014736735139, 
    690.120598847495, 
    531.541303401829, 
    570.540242715219, 
    814.745870899917, 
    717.685672747195, 
    622.944293928841, 
    705.977796061175, 
    756.222787743853, 
    576.764068893996, 
    720.920720355644, 
    755.728806618481, 
    279.48119975364, 
    10.6551346997799, 
    643.214755119168, 
    254.078339088665, 
    810.010243354957, 
    761.689158662835, 
    668.377897435581, 
    702.9617032332, 
    230.784597121318, 
    75.4338647771928, 
    787.015125868431, 
    828.247719844805, 
    906.1499765787, 
    936.401586688516, 
    24.8111522558328, 
    -37.682847104707, 
    -115.671941725165, 
    -269.47263024769, 
    -280.986192590046, 
    -143.506201973687, 
    -122.27327855784, 
    -137.794437651939, 
    -100.020139948385, 
    -195.9763109692, 
    -199.923581410629, 
    -173.747471370461, 
    -228.871809255636, 
    -842.787210556328, 
    -1602.72258210904, 
    -2043.44550454203, 
    -2280.74689998819,
  -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -203.001009878092, 
    -200, 
    -200, 
    -201.784224684268, 
    -239.95569950202, 
    -277.681575106614, 
    -271.4285137074, 
    176.272129112231, 
    497.293451345514, 
    498.642594067274, 
    772.456717479405, 
    297.325124576133, 
    550.42151091641, 
    -77.4165047216266, 
    531.066893672629, 
    658.777626738174, 
    571.271091315943, 
    835.528172637158, 
    881.609001715, 
    657.84663160437, 
    706.167597831564, 
    682.869975091093, 
    682.640490208331, 
    -46.1642507914048, 
    572.485775609034, 
    568.123989630653, 
    622.828662577561, 
    372.890700747154, 
    616.457808200887, 
    1040.3510197365, 
    955.250719965373, 
    758.353563144253, 
    779.631337993489, 
    758.412176484625, 
    671.827988491081, 
    786.788434266776, 
    566.328416839285, 
    386.004923714765, 
    673.816483654607, 
    860.701723626323, 
    484.820343748055, 
    203.494907174102, 
    608.510237750387, 
    662.786705717663, 
    445.823291962247, 
    461.512113718543, 
    82.6118514212072, 
    613.845702133951, 
    506.538514093482, 
    437.74405688107, 
    831.489341462447, 
    367.774456553876, 
    311.336357229898, 
    -20.987707095878, 
    -78.2287265034291, 
    -262.238052237875, 
    -174.473334146906, 
    -139.358442543602, 
    -233.993782692767, 
    -176.204725763166, 
    -249.540493763309, 
    -237.335063340549, 
    -216.728434093857, 
    -432.599629330613, 
    -1419.45848080079, 
    -2006.77979554522, 
    -2267.32669494561, 
    -2427.09662517962,
  -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -276.712791844421, 
    -200, 
    -200, 
    -204.717044902942, 
    -200.404166756659, 
    -245.877095552468, 
    -361.924134885611, 
    -318.354181462681, 
    -158.284136339642, 
    235.664963510776, 
    540.930971912412, 
    817.478366001725, 
    939.396556157949, 
    -15.5775834016299, 
    668.679197065774, 
    434.146933855692, 
    625.702241442638, 
    685.834180654626, 
    904.791868211977, 
    708.984267317036, 
    495.016625181151, 
    894.83293925902, 
    402.875376625527, 
    -178.71459517313, 
    636.706078412952, 
    615.182221774691, 
    370.37841622587, 
    -99.4669481001886, 
    574.194464987897, 
    958.639211127098, 
    973.76232476998, 
    819.242625972324, 
    774.237881744829, 
    750.251248982292, 
    1014.35096661268, 
    859.523353158027, 
    846.330123380211, 
    317.466393751626, 
    815.955884927066, 
    731.459247994926, 
    877.288476121653, 
    581.591735446839, 
    21.4772633464978, 
    558.493200646, 
    663.06590400858, 
    523.578065511228, 
    223.250264630739, 
    147.85205588603, 
    443.800223902652, 
    502.412490977156, 
    746.845077711151, 
    740.914583169866, 
    391.691185638323, 
    56.5026440615024, 
    -86.1925261359722, 
    -162.502108425469, 
    -183.937761253366, 
    -184.293162945002, 
    -144.815111971916, 
    -221.835947250332, 
    -266.638651250858, 
    -306.311837088489, 
    -659.66053462697, 
    -1322.20406284311, 
    -1871.99320011631, 
    -2304.44706464642, 
    -2608.23357576753, 
    -2644.36535729967,
  -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -202.712237779931, 
    -315.722219050663, 
    -382.761565517072, 
    -317.363104456085, 
    -83.1989183148304, 
    579.420136360937, 
    831.479768169948, 
    -88.8097157206041, 
    565.084808823779, 
    838.585862649917, 
    678.308873773552, 
    552.33604936076, 
    527.674540580578, 
    548.554254380219, 
    741.449691123155, 
    787.18340286135, 
    468.112207557952, 
    67.9647829700871, 
    683.001667800165, 
    526.708879165389, 
    304.101842930432, 
    92.5387495164806, 
    626.659612427101, 
    457.777669208174, 
    880.04373654219, 
    932.41355895996, 
    854.095500574398, 
    1046.89628679675, 
    872.19324920586, 
    744.407146389783, 
    727.969719437175, 
    232.27967841841, 
    517.974020126011, 
    638.01819229126, 
    703.339371846745, 
    738.968042345891, 
    400.349948306368, 
    2.24917603873859, 
    439.954314707105, 
    644.5054640818, 
    462.288375337601, 
    60.431409715008, 
    159.536564471339, 
    304.941416117801, 
    419.238311583892, 
    382.972947444252, 
    247.262638869505, 
    193.354736495794, 
    -54.3475914001466, 
    -87.4009428857285, 
    -96.177998177549, 
    -184.461911845447, 
    -133.041586936788, 
    -198.778905804453, 
    -283.598005164512, 
    -372.503393017303, 
    -1301.38131951379, 
    -1829.61693898508, 
    -2334.95508895823, 
    -2577.81369080069, 
    -2660.81516172744, 
    -2750.46330187756,
  -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -201.485843743883, 
    -223.890421375046, 
    -354.711436597389, 
    -405.812513332221, 
    -236.907420281205, 
    -459.591164745917, 
    341.493335734558, 
    513.971458443602, 
    577.180468850812, 
    303.029146841637, 
    569.636529621317, 
    538.61115242252, 
    116.150723954462, 
    397.882687315556, 
    69.0363293233348, 
    98.2401464516772, 
    555.461674407245, 
    337.388507902825, 
    -190.514643245159, 
    213.323893372993, 
    645.986705835569, 
    565.997132842777, 
    744.541899148189, 
    665.207733666905, 
    648.833832837968, 
    828.188479364779, 
    753.983847802848, 
    931.370865440584, 
    441.925592467334, 
    1016.73827689279, 
    134.06168258631, 
    76.7329614669638, 
    893.569606580233, 
    831.250082881023, 
    507.992577521823, 
    398.468018586266, 
    14.8214855855545, 
    196.978572354203, 
    152.598133698017, 
    -11.667265094006, 
    9.47966148925406, 
    1.62549833374251, 
    263.285030441884, 
    525.340084930286, 
    356.932060974303, 
    96.0797723490322, 
    -47.8654620591356, 
    -65.363273322649, 
    -75.0135412152107, 
    -64.1392633378296, 
    -38.9164147782834, 
    -175.682403859206, 
    -259.350183125974, 
    -1055.75527526927, 
    -2148.45834049855, 
    -2558.72968889431, 
    -2699.37733310815, 
    -2696.87977584719, 
    -2717.4638856074, 
    -2654.50499418628,
  -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -210.424058074779, 
    -433.872984195208, 
    -428.785977746979, 
    -176.231996191308, 
    136.466247228599, 
    71.1237123971006, 
    375.047141042031, 
    434.484347921205, 
    570.65294674556, 
    372.634272007231, 
    84.5042969264727, 
    -20.9752012415184, 
    330.141849073554, 
    375.474937251, 
    -26.9630059619264, 
    66.3494318089721, 
    190.263719537359, 
    327.822036230541, 
    816.203149041571, 
    732.915654779418, 
    553.095999936635, 
    550.707526656572, 
    636.431227198114, 
    415.740699802233, 
    424.470215962945, 
    422.29913589801, 
    332.683263054609, 
    371.399733753764, 
    26.2843278824013, 
    -50.4353246910449, 
    128.884437704123, 
    64.2771605452045, 
    74.3112260310756, 
    20.1083307977776, 
    239.832711231536, 
    -13.0923532227547, 
    -98.431423047356, 
    -17.4976454907795, 
    7.16199615447349, 
    64.8025548802496, 
    323.738666773643, 
    375.649587432586, 
    316.514883677878, 
    9.07242948541066, 
    -37.2739035423765, 
    -45.2646189205852, 
    -127.647453387135, 
    -171.48942515191, 
    -556.656286096528, 
    -1349.02660661211, 
    -2425.88018320392, 
    -2943.36336378075, 
    -3218.90837119382, 
    -3275.54269163126, 
    -2660.50930721201, 
    -2593.94488614243, 
    -2308.16669398326,
  -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -246.758762880778, 
    -251.813254498423, 
    -286.774015569745, 
    -453.142171494513, 
    -705.088038830046, 
    -564.327331790739, 
    312.742086724497, 
    9.68219184339865, 
    316.679772277696, 
    478.648727903976, 
    344.457081003391, 
    554.00591521568, 
    421.266921715138, 
    -71.212035085161, 
    792.998763141014, 
    554.250299840327, 
    -74.5217148779752, 
    516.186974665361, 
    442.836665385247, 
    591.069229228515, 
    1016.39384298976, 
    608.58835565498, 
    264.141235605727, 
    907.411732493163, 
    1095.71472865123, 
    734.14368044008, 
    761.993112348364, 
    763.369192783407, 
    617.222905269003, 
    714.112157567492, 
    620.242977872809, 
    601.461220667591, 
    429.190533500246, 
    313.137033353604, 
    44.3383506546857, 
    -67.7765455972179, 
    55.5135394269992, 
    -121.923550321702, 
    24.1974662946864, 
    -19.6204389295013, 
    -102.189105799592, 
    -22.4917682947273, 
    143.797403258682, 
    452.954031513891, 
    240.638120518812, 
    -101.939396364827, 
    -101.047107062174, 
    -97.2364060529025, 
    -694.336402901634, 
    -1558.91453260058, 
    -1213.80825937236, 
    -2448.63007552094, 
    -2661.11202633847, 
    -3190.47119991564, 
    -3493.70138085037, 
    -3680.850683334, 
    -2663.74731113821, 
    -2347.46729708305, 
    -2300,
  -200, 
    -200, 
    -219.933219839184, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -201.965374740481, 
    -200.349929850152, 
    -206.15107249466, 
    -351.109795125031, 
    -637.280621835127, 
    -352.144576893945, 
    -49.4847443485766, 
    105.372091910588, 
    74.4808933812164, 
    215.417283159611, 
    -139.78310256523, 
    -443.439945861716, 
    337.861080951401, 
    71.1523376819187, 
    -112.9486000343, 
    458.548854721083, 
    47.1533669920742, 
    777.275613278593, 
    907.448333449747, 
    595.096352281377, 
    255.771465896897, 
    941.895431877376, 
    1098.49587607731, 
    853.826839075376, 
    834.061556133685, 
    805.776657164297, 
    835.789342147638, 
    675.609012394445, 
    703.786241896608, 
    546.891766461652, 
    545.870523057616, 
    410.341127329417, 
    356.227570088419, 
    18.5174951987223, 
    -102.193160992587, 
    -122.542780803539, 
    -65.7196831911472, 
    -67.099555574905, 
    -125.761908321872, 
    -99.2510461027653, 
    -132.61811631471, 
    -145.549786326337, 
    -121.012454604248, 
    -138.395683352651, 
    -216.415259916605, 
    -578.583840591261, 
    -1882.78365195214, 
    -2430.42617278405, 
    -2713.4092014565, 
    -3116.08877225153, 
    -3417.18663077874, 
    -3966.18061806402, 
    -3913.79244629452, 
    -2740.57904103995, 
    -2378.357712971, 
    -2300, 
    -2300,
  -200, 
    -200, 
    -206.550304827205, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -205.564592993672, 
    -372.504250457008, 
    -406.082524516414, 
    -423.723296119545, 
    -445.832984356169, 
    -477.684076430949, 
    -527.865702877923, 
    -695.542872224919, 
    -764.39902423718, 
    -366.838723072668, 
    -153.113360016232, 
    -55.2022043214271, 
    149.814423574966, 
    148.983577044238, 
    44.2930102505804, 
    363.395944686666, 
    971.785307077922, 
    394.972115729174, 
    1064.51783482465, 
    957.364092913341, 
    886.859055052406, 
    759.740105187908, 
    1023.12777957725, 
    851.223564199213, 
    943.020710559604, 
    835.68445307784, 
    544.280969908092, 
    359.186854453258, 
    247.703230882411, 
    168.468860914565, 
    -13.3590231104641, 
    -111.887614051545, 
    -108.686511269342, 
    -125.73321017386, 
    -127.959167621438, 
    -107.813715315346, 
    -118.495126695408, 
    -109.250636642215, 
    -160.952503697739, 
    -358.201822107888, 
    -1562.81010635226, 
    -1974.16222358528, 
    -2793.12677541908, 
    -3000.74346923829, 
    -3168.78010806845, 
    -3437.15495964982, 
    -3712.95510409742, 
    -3630.04120088341, 
    -2964.92289400689, 
    -2737.29360425377, 
    -2300, 
    -2300, 
    -2300,
  -200, 
    -200, 
    -216.652383180642, 
    -220.38608790245, 
    -231.312167634358, 
    -421.186357752346, 
    -376.846331725596, 
    -206.199596012026, 
    -212.024761524605, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200.353313138477, 
    -252.367586206344, 
    -247.10337956034, 
    -334.127237215282, 
    -501.633380240582, 
    -495.004848680998, 
    -484.539180131934, 
    -592.648911334096, 
    -169.702058563581, 
    -40.0361370618582, 
    3.91973249922951, 
    487.385515911448, 
    491.138616914327, 
    690.469552487571, 
    480.159749969801, 
    278.313052477504, 
    670.783096595411, 
    600.949552324543, 
    496.620458852825, 
    465.276848198164, 
    808.028330282813, 
    788.924958702163, 
    1187.67795197934, 
    1017.87622362503, 
    803.479831323919, 
    450.151677711538, 
    426.614175341566, 
    340.842393084847, 
    378.647441142086, 
    72.5774907296875, 
    -103.23143970686, 
    -101.300746799183, 
    -123.372923838199, 
    -164.604036640882, 
    -163.995929938015, 
    -150.223913334787, 
    -219.057629291591, 
    -1294.20351751659, 
    -2569.53332488776, 
    -2869.98182522731, 
    -2821.47502626631, 
    -3349.61009235105, 
    -3434.64443190555, 
    -3611.08513481593, 
    -3375.74741697578, 
    -3326.36446405391, 
    -2930.88370171318, 
    -2883.72395446024, 
    -2302.65624419038, 
    -2300, 
    -2300, 
    -2300,
  -200, 
    -200, 
    -247.940273586075, 
    -570.653462229493, 
    -327.741577372694, 
    -201.751997517311, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -220.340565616314, 
    -201.062348967036, 
    -149.344594114973, 
    -145.344297367406, 
    -192.64666496439, 
    -354.401789260468, 
    -441.473479592385, 
    -416.45820983767, 
    -447.377521668675, 
    -310.290380646643, 
    -204.363552495055, 
    -68.2772099630036, 
    155.435717179001, 
    414.018513430678, 
    223.395258379148, 
    143.454706118326, 
    233.347471220102, 
    376.015899162671, 
    568.542410966934, 
    519.310034680334, 
    102.962331006139, 
    280.71687697829, 
    1045.49321898901, 
    588.122373378013, 
    646.69165022829, 
    630.92616045569, 
    75.1709410401334, 
    213.373755692103, 
    70.9463121116683, 
    -79.9955454235808, 
    -98.4694175976518, 
    -97.8718264762393, 
    -178.011599097516, 
    -577.025978925666, 
    -631.950933193723, 
    -860.281404775068, 
    -1541.1572958166, 
    -2642.89707015532, 
    -2837.65248283908, 
    -3014.83939329961, 
    -3268.15854647339, 
    -3064.96974310282, 
    -3755.53451667949, 
    -3391.72787598615, 
    -3483.64214793991, 
    -2856.69288835171, 
    -2780.08892579628, 
    -2301.64624378849, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -227.785428663386, 
    -200, 
    -551.910360291453, 
    -248.602883920952, 
    -200.203146123939, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -201.790466148402, 
    -200, 
    -200, 
    -150.675545964771, 
    -152.695929385246, 
    -253.384799728735, 
    -345.347586278284, 
    -377.705000156518, 
    -413.41464206059, 
    -384.99682433074, 
    -299.672907262206, 
    -239.249397662293, 
    -191.689534190523, 
    -93.3396625262549, 
    -72.0838678957805, 
    72.4079121923868, 
    435.312109542445, 
    1036.50661758987, 
    973.409208052108, 
    743.884416586615, 
    1166.74473514538, 
    743.877611551145, 
    247.189351931943, 
    86.3558243272219, 
    -0.939736994234877, 
    335.175713324459, 
    -103.819571479573, 
    -172.400865424524, 
    -155.495133420256, 
    -109.511911821526, 
    -91.0167179865911, 
    -98.0391877495837, 
    -307.208619452019, 
    -2016.7893579874, 
    -2360.09425581265, 
    -2802.18039709351, 
    -2650.936289515, 
    -2925.76573316141, 
    -3033.07895259708, 
    -3211.48680700835, 
    -3076.42756398234, 
    -3810.93647303054, 
    -3954.36182030212, 
    -3556.86603070265, 
    -2660.09551267205, 
    -2420.38983629318, 
    -2309.62283916409, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -345.596859217483, 
    -688.247377197004, 
    -301.185906001187, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -199.72185839731, 
    -176.073922258743, 
    -232.955430574406, 
    -287.930529061517, 
    -322.769973212366, 
    -382.466299473504, 
    -340.085701018671, 
    -279.375458605211, 
    -296.922589160027, 
    -271.001590566433, 
    -233.661162830282, 
    -166.823290123252, 
    -113.992107279224, 
    21.0580688508071, 
    207.478099485537, 
    607.403743363703, 
    714.830351655436, 
    1035.47618967634, 
    774.74440116925, 
    762.519599085829, 
    776.140005720413, 
    241.77793155298, 
    -109.038990467157, 
    -182.886812239988, 
    -676.315953603937, 
    -708.591845581832, 
    -265.385529222314, 
    -237.364286215554, 
    -278.659003246015, 
    -1510.01240577149, 
    -2900.90262657585, 
    -2750.07528221754, 
    -2962.34192844575, 
    -2995.92974327234, 
    -3069.08630063526, 
    -3212.32091171077, 
    -3531.4997554493, 
    -4056.45577452726, 
    -4037.09231987726, 
    -3364.17616823884, 
    -2424.5422783624, 
    -1809.87051649616, 
    -2197.50359601645, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -200.497687515994, 
    -763.214395444043, 
    -218.481519765309, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200.398198968219, 
    -236.483367296245, 
    -200, 
    -200, 
    -200, 
    -202.612320411913, 
    -229.259940167692, 
    -259.094907015196, 
    -286.062966819841, 
    -300.931353937471, 
    -311.308683854601, 
    -307.344404380772, 
    -263.235905486018, 
    -273.192096684574, 
    -269.333430030711, 
    -265.162244999662, 
    -227.545161429873, 
    -177.115417130184, 
    -120.827289556737, 
    -104.556112992136, 
    -65.6389607798535, 
    41.4207558498227, 
    40.9651092879446, 
    103.449890091854, 
    1.83433311569824, 
    27.3187500973866, 
    -104.208058979322, 
    -281.88325294589, 
    -608.672484065767, 
    -1678.20988078188, 
    -2541.03216539067, 
    -2475.09030728915, 
    -1497.59176575942, 
    -2105.7878954846, 
    -2070.850145073, 
    -3097.71954355957, 
    -3018.18232045276, 
    -3169.80556950243, 
    -3201.92134946885, 
    -3315.18512533601, 
    -3894.2560826352, 
    -4471.5804025067, 
    -3997.8971794786, 
    -3222.34974415809, 
    -2365.5919825777, 
    -2338.39802105298, 
    -2304.43890268085, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -344.467311156424, 
    -630.034789949353, 
    -200, 
    -200, 
    -200, 
    -200.164252314295, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200.312523281187, 
    -264.349075610002, 
    -217.451376441879, 
    -200, 
    -200, 
    -200.545078548846, 
    -254.524211872867, 
    -299.383746613849, 
    -304.522848767904, 
    -297.770378685211, 
    -286.510318610863, 
    -295.187657068985, 
    -279.48561664765, 
    -283.073728443928, 
    -293.174736151103, 
    -299.203563536402, 
    -301.72016168148, 
    -292.955082281441, 
    -266.704548680905, 
    -222.780658151643, 
    -174.424698211313, 
    -129.653772234517, 
    -117.065328908795, 
    -127.929949609858, 
    -139.19517114475, 
    -193.782614036212, 
    -207.580424044996, 
    -337.785149530501, 
    -633.14742566118, 
    -1036.99811981988, 
    -1902.44078579996, 
    -2969.59823102621, 
    -3300.18774137252, 
    -2427.36466725382, 
    -2804.95389433003, 
    -3299.65353161171, 
    -3344.65137173267, 
    -3244.59336977763, 
    -3216.97027054773, 
    -3210.33479314208, 
    -4035.71723225458, 
    -4261.37519868889, 
    -3913.51736310078, 
    -2894.61434755397, 
    -2414.45130699986, 
    -2805.24084732382, 
    -3047.08066127387, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -1178.11246650249, 
    -601.134555846554, 
    -200, 
    -203.883904389811, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -228.542060080994, 
    -222.960087140758, 
    -251.999115184599, 
    -206.214685762583, 
    -215.929058102719, 
    -222.300677539788, 
    -280.464623813267, 
    -382.004039277427, 
    -344.964024196682, 
    -302.244164529867, 
    -301.325984412319, 
    -298.288423228504, 
    -281.902633081759, 
    -303.218629155688, 
    -318.492724594852, 
    -327.497771964764, 
    -368.186868174215, 
    -423.75774108443, 
    -486.578514043598, 
    -413.309681545321, 
    -273.056145626382, 
    -196.903352807912, 
    -177.282805764262, 
    -196.284393831705, 
    -207.134306543487, 
    -273.605305743247, 
    -291.968780111761, 
    -850.140009513769, 
    -1739.69918348224, 
    -1931.08423579476, 
    -1996.409370841, 
    -2890.5909576587, 
    -3375.21428172078, 
    -2916.6923056813, 
    -3437.09304098748, 
    -3487.87293201545, 
    -3461.7523216256, 
    -3425.60489824559, 
    -3513.18464802468, 
    -3233.82420463604, 
    -4142.76961559197, 
    -2668.28960368292, 
    -2716.44877619388, 
    -2806.28175068653, 
    -3199.54293047489, 
    -3275.5164424815, 
    -2301.97526562254, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -1822.10257894387, 
    -301.367853391074, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -222.610244415644, 
    -200, 
    -200.158698347888, 
    -207.0966069135, 
    -200, 
    -246.301397379139, 
    -245.016370679336, 
    -219.898779833837, 
    -256.408589928041, 
    -254.600129722349, 
    -334.850593609616, 
    -452.773787307316, 
    -553.485364224052, 
    -469.973071500948, 
    -341.680241775941, 
    -415.025536147374, 
    -333.725261517363, 
    -380.734155964615, 
    -551.356544750959, 
    -739.781279782865, 
    -949.267484111757, 
    -1096.76391762184, 
    -1346.48322192768, 
    -1427.41091701941, 
    -1181.65476422456, 
    -672.235272910549, 
    -363.73214279124, 
    -272.867036595194, 
    -337.037013781168, 
    -498.345810004881, 
    -592.807974906157, 
    -522.71458337663, 
    -633.652264995515, 
    -2828.89529911054, 
    -2340.74227102179, 
    -2023.96552110013, 
    -2936.86661361236, 
    -3465.39463370431, 
    -3491.8772152071, 
    -3092.88439179317, 
    -2885.51023203473, 
    -3864.37629188803, 
    -3852.31645139414, 
    -3528.90805016116, 
    -2844.93968134047, 
    -3137.22510172298, 
    -3155.79646279059, 
    -3753.5018642037, 
    -3994.11488101359, 
    -3486.62597546892, 
    -2331.34695954018, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -1770.72954583248, 
    -219.008961881528, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -206.128297135117, 
    -200, 
    -200, 
    -200, 
    -200, 
    -235.313610835145, 
    -200, 
    -200, 
    -200, 
    -200.131293848941, 
    -220.289754160575, 
    -231.702210850304, 
    -225.262977980286, 
    -254.7570075348, 
    -283.496571774712, 
    -458.420859995775, 
    -598.576305325328, 
    -847.705179417386, 
    -792.186181755108, 
    -757.089620814477, 
    -753.497162941722, 
    -616.42910909279, 
    -1098.79607845875, 
    -1849.00733534246, 
    -2014.2549622163, 
    -1937.67839072506, 
    -1939.10073104124, 
    -2075.97483752209, 
    -2065.19053217598, 
    -1836.08630273697, 
    -1577.76079194516, 
    -848.21635652309, 
    -592.370050120593, 
    -555.557478512789, 
    -796.047147257466, 
    -1030.53594950199, 
    -905.065538446952, 
    -835.835754753361, 
    -2113.81570087703, 
    -1922.58484725696, 
    -2648.17487464213, 
    -3608.637155394, 
    -3593.2795157267, 
    -3643.8395952009, 
    -3443.61130984178, 
    -4015.38112043187, 
    -3927.70928955078, 
    -3566.45749345632, 
    -2683.49924854308, 
    -3251.75598059097, 
    -3551.02076671638, 
    -3996.05143367003, 
    -4368.67428366735, 
    -4149.42346362277, 
    -2518.09102074428, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300 ;
}
