netcdf gmask1m_0 {
dimensions:
	n = 3765 ;
variables:
	int starts(n) ;
	int runlens(n) ;
	int runvals(n) ;
data:

 starts = 
    0, 
    1, 
    2, 
    4, 
    5, 
    10, 
    11, 
    18, 
    19, 
    28, 
    29, 
    40, 
    41, 
    55, 
    56, 
    72, 
    73, 
    91, 
    92, 
    112, 
    113, 
    136, 
    137, 
    163, 
    164, 
    192, 
    193, 
    223, 
    224, 
    257, 
    258, 
    293, 
    294, 
    331, 
    332, 
    371, 
    372, 
    414, 
    415, 
    459, 
    460, 
    506, 
    507, 
    555, 
    556, 
    607, 
    608, 
    661, 
    662, 
    717, 
    718, 
    776, 
    777, 
    837, 
    838, 
    900, 
    901, 
    965, 
    966, 
    1033, 
    1034, 
    1103, 
    1104, 
    1175, 
    1176, 
    1249, 
    1250, 
    1326, 
    1327, 
    1405, 
    1406, 
    1486, 
    1487, 
    1569, 
    1570, 
    1655, 
    1656, 
    1743, 
    1744, 
    1833, 
    1834, 
    1925, 
    1926, 
    2021, 
    2022, 
    2119, 
    2120, 
    2219, 
    2220, 
    2321, 
    2322, 
    2426, 
    2427, 
    2533, 
    2534, 
    2642, 
    2643, 
    2753, 
    2754, 
    2867, 
    2868, 
    2983, 
    2984, 
    3101, 
    3102, 
    3222, 
    3223, 
    3345, 
    3346, 
    3470, 
    3471, 
    3597, 
    3598, 
    3727, 
    3728, 
    3859, 
    3860, 
    3993, 
    3994, 
    4129, 
    4130, 
    4268, 
    4269, 
    4409, 
    4410, 
    4552, 
    4553, 
    4697, 
    4698, 
    4845, 
    4846, 
    4995, 
    4996, 
    5147, 
    5148, 
    5301, 
    5302, 
    5458, 
    5459, 
    5617, 
    5618, 
    5778, 
    5779, 
    5942, 
    5943, 
    6109, 
    6110, 
    6278, 
    6279, 
    6449, 
    6450, 
    6623, 
    6624, 
    6799, 
    6800, 
    6977, 
    6978, 
    7157, 
    7158, 
    7340, 
    7341, 
    7525, 
    7526, 
    7712, 
    7713, 
    7901, 
    7902, 
    8093, 
    8094, 
    8287, 
    8288, 
    8483, 
    8484, 
    8681, 
    8682, 
    8882, 
    8883, 
    9085, 
    9086, 
    9290, 
    9291, 
    9497, 
    9498, 
    9707, 
    9708, 
    9919, 
    9920, 
    10133, 
    10134, 
    10349, 
    10350, 
    10568, 
    10569, 
    10789, 
    10790, 
    11012, 
    11013, 
    11237, 
    11238, 
    11465, 
    11466, 
    11695, 
    11696, 
    11927, 
    11928, 
    12163, 
    12164, 
    12401, 
    12402, 
    12641, 
    12642, 
    12883, 
    12884, 
    13128, 
    13129, 
    13375, 
    13376, 
    13624, 
    13625, 
    13875, 
    13876, 
    14129, 
    14130, 
    14385, 
    14386, 
    14643, 
    14644, 
    14903, 
    14904, 
    15166, 
    15167, 
    15431, 
    15432, 
    15698, 
    15699, 
    15967, 
    15968, 
    16239, 
    16240, 
    16513, 
    16514, 
    16789, 
    16790, 
    17067, 
    17068, 
    17348, 
    17349, 
    17631, 
    17632, 
    17916, 
    17917, 
    18204, 
    18205, 
    18494, 
    18495, 
    18786, 
    18787, 
    19080, 
    19081, 
    19377, 
    19378, 
    19676, 
    19677, 
    19977, 
    19978, 
    20281, 
    20282, 
    20588, 
    20589, 
    20897, 
    20898, 
    21208, 
    21209, 
    21521, 
    21522, 
    21837, 
    21838, 
    22155, 
    22156, 
    22475, 
    22476, 
    22797, 
    22798, 
    23122, 
    23123, 
    23449, 
    23450, 
    23778, 
    23779, 
    24109, 
    24110, 
    24443, 
    24444, 
    24779, 
    24780, 
    25117, 
    25118, 
    25457, 
    25458, 
    25800, 
    25801, 
    26145, 
    26146, 
    26492, 
    26493, 
    26842, 
    26843, 
    27194, 
    27195, 
    27548, 
    27549, 
    27904, 
    27905, 
    28263, 
    28264, 
    28624, 
    28625, 
    28987, 
    28988, 
    29352, 
    29353, 
    29720, 
    29721, 
    30090, 
    30091, 
    30462, 
    30463, 
    30837, 
    30838, 
    31215, 
    31216, 
    31595, 
    31596, 
    31977, 
    31978, 
    32361, 
    32362, 
    32748, 
    32749, 
    33137, 
    33138, 
    33528, 
    33529, 
    33921, 
    33922, 
    34317, 
    34318, 
    34715, 
    34716, 
    35115, 
    35116, 
    35518, 
    35519, 
    35923, 
    35924, 
    36330, 
    36331, 
    36739, 
    36740, 
    37151, 
    37152, 
    37565, 
    37566, 
    37981, 
    37982, 
    38399, 
    38400, 
    38820, 
    38821, 
    39243, 
    39244, 
    39668, 
    39669, 
    40095, 
    40096, 
    40525, 
    40526, 
    40957, 
    40958, 
    41391, 
    41392, 
    41827, 
    41828, 
    42266, 
    42267, 
    42707, 
    42708, 
    43151, 
    43152, 
    43597, 
    43598, 
    44046, 
    44047, 
    44497, 
    44498, 
    44950, 
    44951, 
    45405, 
    45406, 
    45863, 
    45864, 
    46323, 
    46324, 
    46785, 
    46786, 
    47250, 
    47251, 
    47717, 
    47718, 
    48186, 
    48187, 
    48657, 
    48658, 
    49131, 
    49132, 
    49607, 
    49608, 
    50085, 
    50086, 
    50565, 
    50566, 
    51048, 
    51049, 
    51533, 
    51534, 
    52020, 
    52021, 
    52509, 
    52510, 
    53001, 
    53002, 
    53495, 
    53496, 
    53991, 
    53992, 
    54489, 
    54490, 
    54990, 
    54991, 
    55493, 
    55494, 
    55998, 
    55999, 
    56505, 
    56506, 
    57015, 
    57016, 
    57528, 
    57529, 
    58043, 
    58044, 
    58561, 
    58562, 
    59081, 
    59082, 
    59603, 
    59604, 
    60127, 
    60128, 
    60654, 
    60655, 
    61183, 
    61184, 
    61714, 
    61715, 
    62247, 
    62248, 
    62783, 
    62784, 
    63321, 
    63322, 
    63861, 
    63862, 
    64403, 
    64404, 
    64948, 
    64949, 
    65495, 
    65496, 
    66044, 
    66045, 
    66595, 
    66596, 
    67149, 
    67150, 
    67705, 
    67706, 
    68263, 
    68264, 
    68823, 
    68824, 
    69386, 
    69387, 
    69951, 
    69952, 
    70518, 
    70519, 
    71087, 
    71088, 
    71659, 
    71660, 
    72233, 
    72234, 
    72809, 
    72810, 
    73388, 
    73389, 
    73970, 
    73971, 
    74554, 
    74555, 
    75140, 
    75141, 
    75729, 
    75730, 
    76320, 
    76321, 
    76913, 
    76914, 
    77508, 
    77509, 
    78106, 
    78107, 
    78706, 
    78707, 
    79308, 
    79309, 
    79912, 
    79913, 
    80519, 
    80520, 
    81128, 
    81129, 
    81739, 
    81740, 
    82352, 
    82353, 
    82968, 
    82969, 
    83586, 
    83587, 
    84206, 
    84207, 
    84828, 
    84829, 
    85453, 
    85454, 
    86080, 
    86081, 
    86709, 
    86710, 
    87341, 
    87342, 
    87975, 
    87976, 
    88611, 
    88612, 
    89249, 
    89250, 
    89890, 
    89891, 
    90533, 
    90534, 
    91178, 
    91179, 
    91825, 
    91826, 
    92475, 
    92476, 
    93128, 
    93129, 
    93783, 
    93784, 
    94440, 
    94441, 
    95100, 
    95101, 
    95762, 
    95763, 
    96426, 
    96427, 
    97092, 
    97093, 
    97761, 
    97762, 
    98432, 
    98433, 
    99105, 
    99106, 
    99780, 
    99781, 
    100458, 
    100459, 
    101138, 
    101139, 
    101820, 
    101821, 
    102504, 
    102505, 
    103191, 
    103192, 
    103880, 
    103881, 
    104571, 
    104572, 
    105265, 
    105266, 
    105961, 
    105962, 
    106659, 
    106660, 
    107359, 
    107360, 
    108062, 
    108063, 
    108767, 
    108768, 
    109474, 
    109475, 
    110183, 
    110184, 
    110895, 
    110896, 
    111609, 
    111610, 
    112325, 
    112326, 
    113043, 
    113044, 
    113764, 
    113765, 
    114488, 
    114489, 
    115214, 
    115215, 
    115942, 
    115943, 
    116673, 
    116674, 
    117406, 
    117407, 
    118141, 
    118142, 
    118878, 
    118879, 
    119618, 
    119619, 
    120360, 
    120361, 
    121104, 
    121105, 
    121851, 
    121852, 
    122600, 
    122601, 
    123351, 
    123352, 
    124104, 
    124105, 
    124860, 
    124861, 
    125618, 
    125619, 
    126378, 
    126379, 
    127140, 
    127141, 
    127905, 
    127906, 
    128672, 
    128673, 
    129441, 
    129442, 
    130212, 
    130213, 
    130986, 
    130987, 
    131762, 
    131763, 
    132540, 
    132541, 
    133320, 
    133321, 
    134103, 
    134104, 
    134888, 
    134889, 
    135675, 
    135676, 
    136464, 
    136465, 
    137257, 
    137258, 
    138052, 
    138053, 
    138849, 
    138850, 
    139648, 
    139649, 
    140450, 
    140451, 
    141254, 
    141255, 
    142060, 
    142061, 
    142869, 
    142870, 
    143680, 
    143681, 
    144493, 
    144494, 
    145308, 
    145309, 
    146126, 
    146127, 
    146946, 
    146947, 
    147768, 
    147769, 
    148592, 
    148593, 
    149419, 
    149420, 
    150248, 
    150249, 
    151079, 
    151080, 
    151912, 
    151913, 
    152748, 
    152749, 
    153586, 
    153587, 
    154426, 
    154427, 
    155268, 
    155269, 
    156113, 
    156114, 
    156960, 
    156961, 
    157809, 
    157810, 
    158660, 
    158661, 
    159514, 
    159515, 
    160370, 
    160371, 
    161228, 
    161229, 
    162090, 
    162091, 
    162954, 
    162955, 
    163820, 
    163821, 
    164688, 
    164689, 
    165559, 
    165560, 
    166432, 
    166433, 
    167307, 
    167308, 
    168184, 
    168185, 
    169064, 
    169065, 
    169946, 
    169947, 
    170830, 
    170831, 
    171716, 
    171717, 
    172605, 
    172606, 
    173496, 
    173497, 
    174389, 
    174390, 
    175284, 
    175285, 
    176182, 
    176183, 
    177082, 
    177083, 
    177984, 
    177985, 
    178888, 
    178889, 
    179795, 
    179796, 
    180704, 
    180705, 
    181615, 
    181616, 
    182528, 
    182529, 
    183444, 
    183445, 
    184362, 
    184363, 
    185282, 
    185283, 
    186204, 
    186205, 
    187129, 
    187130, 
    188056, 
    188057, 
    188985, 
    188986, 
    189918, 
    189919, 
    190853, 
    190854, 
    191790, 
    191791, 
    192729, 
    192730, 
    193671, 
    193672, 
    194615, 
    194616, 
    195561, 
    195562, 
    196509, 
    196510, 
    197460, 
    197461, 
    198413, 
    198414, 
    199368, 
    199369, 
    200325, 
    200326, 
    201285, 
    201286, 
    202247, 
    202248, 
    203211, 
    203212, 
    204177, 
    204178, 
    205146, 
    205147, 
    206117, 
    206118, 
    207090, 
    207091, 
    208066, 
    208067, 
    209044, 
    209045, 
    210024, 
    210025, 
    211006, 
    211007, 
    211991, 
    211992, 
    212978, 
    212979, 
    213967, 
    213968, 
    214958, 
    214959, 
    215952, 
    215953, 
    216948, 
    216949, 
    217946, 
    217947, 
    218947, 
    218948, 
    219951, 
    219952, 
    220957, 
    220958, 
    221965, 
    221966, 
    222975, 
    222976, 
    223988, 
    223989, 
    225003, 
    225004, 
    226020, 
    226021, 
    227039, 
    227040, 
    228061, 
    228062, 
    229085, 
    229086, 
    230111, 
    230112, 
    231139, 
    231140, 
    232170, 
    232171, 
    233203, 
    233204, 
    234238, 
    234239, 
    235275, 
    235276, 
    236315, 
    236316, 
    237357, 
    237358, 
    238401, 
    238402, 
    239448, 
    239449, 
    240497, 
    240498, 
    241548, 
    241549, 
    242601, 
    242602, 
    243657, 
    243658, 
    244715, 
    244716, 
    245775, 
    245776, 
    246837, 
    246838, 
    247902, 
    247903, 
    248969, 
    248970, 
    250038, 
    250039, 
    251110, 
    251111, 
    252185, 
    252186, 
    253262, 
    253263, 
    254341, 
    254342, 
    255422, 
    255423, 
    256506, 
    256507, 
    257592, 
    257593, 
    258680, 
    258681, 
    259771, 
    259772, 
    260864, 
    260865, 
    261959, 
    261960, 
    263056, 
    263057, 
    264156, 
    264157, 
    265258, 
    265259, 
    266362, 
    266363, 
    267468, 
    267469, 
    268577, 
    268578, 
    269688, 
    269689, 
    270801, 
    270802, 
    271916, 
    271917, 
    273034, 
    273035, 
    274154, 
    274155, 
    275276, 
    275277, 
    276400, 
    276401, 
    277527, 
    277528, 
    278656, 
    278657, 
    279787, 
    279788, 
    280920, 
    280921, 
    282056, 
    282057, 
    283194, 
    283195, 
    284335, 
    284336, 
    285478, 
    285479, 
    286624, 
    286625, 
    287772, 
    287773, 
    288922, 
    288923, 
    290075, 
    290076, 
    291230, 
    291231, 
    292387, 
    292388, 
    293546, 
    293547, 
    294708, 
    294709, 
    295872, 
    295873, 
    297038, 
    297039, 
    298206, 
    298207, 
    299377, 
    299378, 
    300550, 
    300551, 
    301725, 
    301726, 
    302902, 
    302903, 
    304082, 
    304083, 
    305264, 
    305265, 
    306448, 
    306449, 
    307634, 
    307635, 
    308823, 
    308824, 
    310014, 
    310015, 
    311207, 
    311208, 
    312402, 
    312403, 
    313600, 
    313601, 
    314800, 
    314801, 
    316002, 
    316003, 
    317207, 
    317208, 
    318414, 
    318415, 
    319624, 
    319625, 
    320836, 
    320837, 
    322051, 
    322052, 
    323268, 
    323269, 
    324487, 
    324488, 
    325708, 
    325709, 
    326932, 
    326933, 
    328158, 
    328159, 
    329386, 
    329387, 
    330616, 
    330617, 
    331849, 
    331850, 
    333084, 
    333085, 
    334321, 
    334322, 
    335560, 
    335561, 
    336802, 
    336803, 
    338046, 
    338047, 
    339292, 
    339293, 
    340540, 
    340541, 
    341791, 
    341792, 
    343044, 
    343045, 
    344299, 
    344300, 
    345556, 
    345557, 
    346816, 
    346817, 
    348078, 
    348079, 
    349342, 
    349343, 
    350609, 
    350610, 
    351878, 
    351879, 
    353149, 
    353150, 
    354422, 
    354423, 
    355698, 
    355699, 
    356976, 
    356977, 
    358257, 
    358258, 
    359540, 
    359541, 
    360826, 
    360827, 
    362114, 
    362115, 
    363404, 
    363405, 
    364696, 
    364697, 
    365991, 
    365992, 
    367288, 
    367289, 
    368587, 
    368588, 
    369888, 
    369889, 
    371192, 
    371193, 
    372498, 
    372499, 
    373806, 
    373807, 
    375116, 
    375117, 
    376429, 
    376430, 
    377744, 
    377745, 
    379061, 
    379062, 
    380381, 
    380382, 
    381703, 
    381704, 
    383027, 
    383028, 
    384353, 
    384354, 
    385682, 
    385683, 
    387013, 
    387014, 
    388346, 
    388347, 
    389681, 
    389682, 
    391019, 
    391020, 
    392359, 
    392360, 
    393701, 
    393702, 
    395045, 
    395046, 
    396392, 
    396393, 
    397742, 
    397743, 
    399094, 
    399095, 
    400448, 
    400449, 
    401805, 
    401806, 
    403164, 
    403165, 
    404525, 
    404526, 
    405888, 
    405889, 
    407254, 
    407255, 
    408622, 
    408623, 
    409992, 
    409993, 
    411364, 
    411365, 
    412739, 
    412740, 
    414116, 
    414117, 
    415495, 
    415496, 
    416877, 
    416878, 
    418261, 
    418262, 
    419647, 
    419648, 
    421035, 
    421036, 
    422426, 
    422427, 
    423819, 
    423820, 
    425214, 
    425215, 
    426611, 
    426612, 
    428011, 
    428012, 
    429413, 
    429414, 
    430817, 
    430818, 
    432223, 
    432224, 
    433632, 
    433633, 
    435043, 
    435044, 
    436456, 
    436457, 
    437871, 
    437872, 
    439289, 
    439290, 
    440710, 
    440711, 
    442133, 
    442134, 
    443558, 
    443559, 
    444986, 
    444987, 
    446416, 
    446417, 
    447848, 
    447849, 
    449283, 
    449284, 
    450720, 
    450721, 
    452159, 
    452160, 
    453600, 
    453601, 
    455044, 
    455045, 
    456490, 
    456491, 
    457938, 
    457939, 
    459388, 
    459389, 
    460841, 
    460842, 
    462296, 
    462297, 
    463753, 
    463754, 
    465212, 
    465213, 
    466674, 
    466675, 
    468138, 
    468139, 
    469604, 
    469605, 
    471072, 
    471073, 
    472543, 
    472544, 
    474016, 
    474017, 
    475491, 
    475492, 
    476968, 
    476969, 
    478448, 
    478449, 
    479930, 
    479931, 
    481414, 
    481415, 
    482900, 
    482901, 
    484390, 
    484391, 
    485882, 
    485883, 
    487376, 
    487377, 
    488873, 
    488874, 
    490372, 
    490373, 
    491873, 
    491874, 
    493376, 
    493377, 
    494882, 
    494883, 
    496390, 
    496391, 
    497900, 
    497901, 
    499412, 
    499413, 
    500927, 
    500928, 
    502444, 
    502445, 
    503963, 
    503964, 
    505484, 
    505485, 
    507008, 
    507009, 
    508534, 
    508535, 
    510062, 
    510063, 
    511594, 
    511595, 
    513131, 
    513132, 
    514673, 
    514674, 
    516219, 
    516220, 
    517770, 
    517771, 
    519325, 
    519326, 
    520885, 
    520886, 
    522449, 
    522450, 
    524018, 
    524019, 
    525592, 
    525593, 
    527170, 
    527171, 
    528753, 
    528754, 
    530341, 
    530342, 
    531934, 
    531935, 
    533531, 
    533532, 
    535133, 
    535134, 
    536740, 
    536741, 
    538351, 
    538352, 
    539967, 
    539968, 
    541587, 
    541588, 
    543212, 
    543213, 
    544841, 
    544842, 
    546475, 
    546476, 
    548113, 
    548114, 
    549756, 
    549757, 
    551404, 
    551405, 
    553056, 
    553057, 
    554713, 
    554714, 
    556374, 
    556375, 
    558040, 
    558041, 
    559710, 
    559711, 
    561385, 
    561386, 
    563065, 
    563066, 
    564749, 
    564750, 
    566438, 
    566439, 
    568131, 
    568132, 
    569829, 
    569830, 
    571531, 
    571532, 
    573238, 
    573239, 
    574950, 
    574951, 
    576666, 
    576667, 
    578387, 
    578388, 
    580112, 
    580113, 
    581843, 
    581844, 
    583578, 
    583579, 
    585318, 
    585319, 
    587063, 
    587064, 
    588812, 
    588813, 
    590566, 
    590567, 
    592324, 
    592325, 
    594087, 
    594088, 
    595854, 
    595855, 
    597626, 
    597627, 
    599402, 
    599403, 
    601183, 
    601184, 
    602969, 
    602970, 
    604759, 
    604760, 
    606554, 
    606555, 
    608353, 
    608354, 
    610157, 
    610158, 
    611965, 
    611966, 
    613778, 
    613779, 
    615596, 
    615597, 
    617418, 
    617419, 
    619245, 
    619246, 
    621076, 
    621077, 
    622912, 
    622913, 
    624752, 
    624753, 
    626597, 
    626598, 
    628447, 
    628448, 
    630301, 
    630302, 
    632160, 
    632161, 
    634023, 
    634024, 
    635892, 
    635893, 
    637765, 
    637766, 
    639643, 
    639644, 
    641526, 
    641527, 
    643413, 
    643414, 
    645305, 
    645306, 
    647201, 
    647202, 
    649102, 
    649103, 
    651007, 
    651008, 
    652917, 
    652918, 
    654831, 
    654832, 
    656750, 
    656751, 
    658673, 
    658674, 
    660601, 
    660602, 
    662534, 
    662535, 
    664471, 
    664472, 
    666413, 
    666414, 
    668359, 
    668360, 
    670310, 
    670311, 
    672266, 
    672267, 
    674226, 
    674227, 
    676191, 
    676192, 
    678160, 
    678161, 
    680134, 
    680135, 
    682112, 
    682113, 
    684095, 
    684096, 
    686083, 
    686084, 
    688075, 
    688076, 
    690072, 
    690073, 
    692073, 
    692074, 
    694079, 
    694080, 
    696090, 
    696091, 
    698106, 
    698107, 
    700127, 
    700128, 
    702152, 
    702153, 
    704182, 
    704183, 
    706216, 
    706217, 
    708255, 
    708256, 
    710298, 
    710299, 
    712346, 
    712347, 
    714398, 
    714399, 
    716455, 
    716456, 
    718517, 
    718518, 
    720583, 
    720584, 
    722654, 
    722655, 
    724729, 
    724730, 
    726809, 
    726810, 
    728893, 
    728894, 
    730982, 
    730983, 
    733076, 
    733077, 
    735174, 
    735175, 
    737277, 
    737278, 
    739384, 
    739385, 
    741496, 
    741497, 
    743612, 
    743613, 
    745733, 
    745734, 
    747859, 
    747860, 
    749989, 
    749990, 
    752124, 
    752125, 
    754263, 
    754264, 
    756407, 
    756408, 
    758556, 
    758557, 
    760710, 
    760711, 
    762869, 
    762870, 
    765032, 
    765033, 
    767200, 
    767201, 
    769372, 
    769373, 
    771549, 
    771550, 
    773730, 
    773731, 
    775916, 
    775917, 
    778106, 
    778107, 
    780301, 
    780302, 
    782501, 
    782502, 
    784705, 
    784706, 
    786914, 
    786915, 
    789127, 
    789128, 
    791345, 
    791346, 
    793567, 
    793568, 
    795794, 
    795795, 
    798026, 
    798027, 
    800262, 
    800263, 
    802503, 
    802504, 
    804748, 
    804749, 
    806998, 
    806999, 
    809252, 
    809253, 
    811511, 
    811512, 
    813775, 
    813776, 
    816043, 
    816044, 
    818316, 
    818317, 
    820593, 
    820594, 
    822875, 
    822876, 
    825162, 
    825163, 
    827454, 
    827455, 
    829751, 
    829752, 
    832052, 
    832053, 
    834358, 
    834359, 
    836668, 
    836669, 
    838983, 
    838984, 
    841302, 
    841303, 
    843626, 
    843627, 
    845954, 
    845955, 
    848287, 
    848288, 
    850624, 
    850625, 
    852966, 
    852967, 
    855313, 
    855314, 
    857664, 
    857665, 
    860020, 
    860021, 
    862380, 
    862381, 
    864745, 
    864746, 
    867115, 
    867116, 
    869489, 
    869490, 
    871868, 
    871869, 
    874251, 
    874252, 
    876639, 
    876640, 
    879031, 
    879032, 
    881428, 
    881429, 
    883830, 
    883831, 
    886236, 
    886237, 
    888647, 
    888648, 
    891062, 
    891063, 
    893482, 
    893483, 
    895906, 
    895907, 
    898336, 
    898337, 
    900771, 
    900772, 
    903210, 
    903211, 
    905654, 
    905655, 
    908102, 
    908103, 
    910552, 
    910553, 
    913004, 
    913005, 
    915458, 
    915459, 
    917913, 
    917914, 
    920370, 
    920371, 
    922829, 
    922830, 
    925289, 
    925290, 
    927751, 
    927752, 
    930215, 
    930216, 
    932681, 
    932682, 
    935148, 
    935149, 
    937617, 
    937618, 
    940088, 
    940089, 
    942560, 
    942561, 
    945034, 
    945035, 
    947510, 
    947511, 
    949987, 
    949988, 
    952466, 
    952467, 
    954947, 
    954948, 
    957430, 
    957431, 
    959914, 
    959915, 
    962400, 
    962401, 
    964888, 
    964889, 
    967377, 
    967378, 
    969868, 
    969869, 
    972362, 
    972363, 
    974857, 
    974858, 
    977354, 
    977355, 
    979853, 
    979854, 
    982354, 
    982355, 
    984856, 
    984857, 
    987360, 
    987361, 
    989866, 
    989867, 
    992373, 
    992374, 
    994882, 
    994883, 
    997393, 
    997394, 
    999905, 
    999906, 
    1002419, 
    1002420, 
    1004935, 
    1004936, 
    1007453, 
    1007454, 
    1009972, 
    1009973, 
    1012493, 
    1012494, 
    1015016, 
    1015017, 
    1017540, 
    1017541, 
    1020066, 
    1020067, 
    1022594, 
    1022595, 
    1025123, 
    1025124, 
    1027654, 
    1027655, 
    1030187, 
    1030188, 
    1032722, 
    1032723, 
    1035258, 
    1035259, 
    1037796, 
    1037797, 
    1040336, 
    1040337, 
    1042877, 
    1042878, 
    1045420, 
    1045421, 
    1047965, 
    1047966, 
    1050512, 
    1050513, 
    1053061, 
    1053062, 
    1055612, 
    1055613, 
    1058165, 
    1058166, 
    1060719, 
    1060720, 
    1063275, 
    1063276, 
    1065833, 
    1065834, 
    1068392, 
    1068393, 
    1070953, 
    1070954, 
    1073516, 
    1073517, 
    1076080, 
    1076081, 
    1078646, 
    1078647, 
    1081214, 
    1081215, 
    1083784, 
    1083785, 
    1086355, 
    1086356, 
    1088928, 
    1088929, 
    1091503, 
    1091504, 
    1094079, 
    1094080, 
    1096657, 
    1096658, 
    1099237, 
    1099238, 
    1101818, 
    1101819, 
    1104401, 
    1104402, 
    1106986, 
    1106987, 
    1109573, 
    1109574, 
    1112161, 
    1112162, 
    1114751, 
    1114752, 
    1117343, 
    1117344, 
    1119936, 
    1119937, 
    1122531, 
    1122532, 
    1125128, 
    1125129, 
    1127727, 
    1127728, 
    1130328, 
    1130329, 
    1132931, 
    1132932, 
    1135536, 
    1135537, 
    1138142, 
    1138143, 
    1140750, 
    1140751, 
    1143360, 
    1143361, 
    1145971, 
    1145972, 
    1148584, 
    1148585, 
    1151199, 
    1151200, 
    1153815, 
    1153816, 
    1156433, 
    1156434, 
    1159053, 
    1159054, 
    1161674, 
    1161675, 
    1164297, 
    1164298, 
    1166922, 
    1166923, 
    1169549, 
    1169550, 
    1172177, 
    1172178, 
    1174807, 
    1174808, 
    1177439, 
    1177440, 
    1180072, 
    1180073, 
    1182707, 
    1182708, 
    1185344, 
    1185345, 
    1187982, 
    1187983, 
    1190622, 
    1190623, 
    1193264, 
    1193265, 
    1195908, 
    1195909, 
    1198553, 
    1198554, 
    1201200, 
    1201201, 
    1203849, 
    1203850, 
    1206500, 
    1206501, 
    1209153, 
    1209154, 
    1211808, 
    1211809, 
    1214464, 
    1214465, 
    1217122, 
    1217123, 
    1219782, 
    1219783, 
    1222444, 
    1222445, 
    1225107, 
    1225108, 
    1227772, 
    1227773, 
    1230439, 
    1230440, 
    1233107, 
    1233108, 
    1235777, 
    1235778, 
    1238449, 
    1238450, 
    1241122, 
    1241123, 
    1243797, 
    1243798, 
    1246474, 
    1246475, 
    1249153, 
    1249154, 
    1251833, 
    1251834, 
    1254515, 
    1254516, 
    1257199, 
    1257200, 
    1259884, 
    1259885, 
    1262571, 
    1262572, 
    1265260, 
    1265261, 
    1267950, 
    1267951, 
    1270642, 
    1270643, 
    1273336, 
    1273337, 
    1276032, 
    1276033, 
    1278729, 
    1278730, 
    1281428, 
    1281429, 
    1284129, 
    1284130, 
    1286832, 
    1286833, 
    1289539, 
    1289540, 
    1292249, 
    1292250, 
    1294962, 
    1294963, 
    1297679, 
    1297680, 
    1300400, 
    1300401, 
    1303125, 
    1303126, 
    1305852, 
    1305853, 
    1308583, 
    1308584, 
    1311318, 
    1311319, 
    1314056, 
    1314057, 
    1316798, 
    1316799, 
    1319543, 
    1319544, 
    1322291, 
    1322292, 
    1325043, 
    1325044, 
    1327799, 
    1327800, 
    1330559, 
    1330560, 
    1333321, 
    1333322, 
    1336087, 
    1336088, 
    1338857, 
    1338858, 
    1341630, 
    1341631, 
    1344407, 
    1344408, 
    1347187, 
    1347188, 
    1349970, 
    1349971, 
    1352757, 
    1352758, 
    1355548, 
    1355549, 
    1358342, 
    1358343, 
    1361139, 
    1361140, 
    1363940, 
    1363941, 
    1366745, 
    1366746, 
    1369553, 
    1369554, 
    1372364, 
    1372365, 
    1375179, 
    1375180, 
    1377997, 
    1377998, 
    1380819, 
    1380820, 
    1383645, 
    1383646, 
    1386474, 
    1386475, 
    1389306, 
    1389307, 
    1392142, 
    1392143, 
    1394982, 
    1394983, 
    1397825, 
    1397826, 
    1400671, 
    1400672, 
    1403521, 
    1403522, 
    1406374, 
    1406375, 
    1409231, 
    1409232, 
    1412092, 
    1412093, 
    1414956, 
    1414957, 
    1417823, 
    1417824, 
    1420694, 
    1420695, 
    1423569, 
    1423570, 
    1426447, 
    1426448, 
    1429328, 
    1429329, 
    1432213, 
    1432214, 
    1435101, 
    1435102, 
    1437993, 
    1437994, 
    1440889, 
    1440890, 
    1443788, 
    1443789, 
    1446690, 
    1446691, 
    1449596, 
    1449597, 
    1452506, 
    1452507, 
    1455419, 
    1455420, 
    1458335, 
    1458336, 
    1461255, 
    1461256, 
    1464178, 
    1464179, 
    1467105, 
    1467106, 
    1470036, 
    1470037, 
    1472970, 
    1472971, 
    1475907, 
    1475908, 
    1478848, 
    1478849, 
    1481793, 
    1481794, 
    1484741, 
    1484742, 
    1487692, 
    1487693, 
    1490647, 
    1490648, 
    1493605, 
    1493606, 
    1496567, 
    1496568, 
    1499533, 
    1499534, 
    1502502, 
    1502503, 
    1505474, 
    1505475, 
    1508450, 
    1508451, 
    1511430, 
    1511431, 
    1514413, 
    1514414, 
    1517399, 
    1517400, 
    1520389, 
    1520390, 
    1523382, 
    1523383, 
    1526379, 
    1526380, 
    1529380, 
    1529381, 
    1532384, 
    1532385, 
    1535391, 
    1535392, 
    1538402, 
    1538403, 
    1541417, 
    1541418, 
    1544435, 
    1544436, 
    1547456, 
    1547457, 
    1550481, 
    1550482, 
    1553509, 
    1553510, 
    1556541, 
    1556542, 
    1559576, 
    1559577, 
    1562615, 
    1562616, 
    1565657, 
    1565658, 
    1568703, 
    1568704, 
    1571753, 
    1571754, 
    1574805, 
    1574806, 
    1577861, 
    1577862, 
    1580921, 
    1580922, 
    1583984, 
    1583985, 
    1587051, 
    1587052, 
    1590121, 
    1590122, 
    1593195, 
    1593196, 
    1596272, 
    1596273, 
    1599353, 
    1599354, 
    1602438, 
    1602439, 
    1605525, 
    1605526, 
    1608616, 
    1608617, 
    1611711, 
    1611712, 
    1614809, 
    1614810, 
    1617911, 
    1617912, 
    1621016, 
    1621017, 
    1624125, 
    1624126, 
    1627237, 
    1627238, 
    1630353, 
    1630354, 
    1633473, 
    1633474, 
    1636595, 
    1636596, 
    1639721, 
    1639722, 
    1642851, 
    1642852, 
    1645984, 
    1645985, 
    1649121, 
    1649122, 
    1652261, 
    1652262, 
    1655405, 
    1655406, 
    1658552, 
    1658553, 
    1661703, 
    1661704, 
    1664858, 
    1664859, 
    1668015, 
    1668016, 
    1671176, 
    1671177, 
    1674341, 
    1674342, 
    1677509, 
    1677510, 
    1680681, 
    1680682, 
    1683856, 
    1683857, 
    1687035, 
    1687036, 
    1690217, 
    1690218, 
    1693403, 
    1693404, 
    1696593, 
    1696594, 
    1699785, 
    1699786, 
    1702981, 
    1702982, 
    1706181, 
    1706182, 
    1709384, 
    1709385, 
    1712591, 
    1712592, 
    1715801, 
    1715802, 
    1719015, 
    1719016, 
    1722232, 
    1722233, 
    1725453, 
    1725454, 
    1728678, 
    1728679, 
    1731905, 
    1731906, 
    1735136, 
    1735137, 
    1738371, 
    1738372, 
    1741609, 
    1741610, 
    1744851, 
    1744852, 
    1748096, 
    1748097, 
    1751345, 
    1751346, 
    1754597, 
    1754598, 
    1757853, 
    1757854, 
    1761113, 
    1761114, 
    1764375, 
    1764376, 
    1767641, 
    1767642, 
    1770911, 
    1770912, 
    1774184, 
    1774185, 
    1777460, 
    1777461, 
    1780740, 
    1780741, 
    1784023, 
    1784024, 
    1787310, 
    1787311, 
    1790601, 
    1790602, 
    1793895, 
    1793896, 
    1797192, 
    1797193, 
    1800493, 
    1800494, 
    1803798, 
    1803799, 
    1807106, 
    1807107, 
    1810417, 
    1810418, 
    1813732, 
    1813733, 
    1817050, 
    1817051, 
    1820372, 
    1820373, 
    1823698, 
    1823699, 
    1827027, 
    1827028, 
    1830359, 
    1830360, 
    1833695, 
    1833696, 
    1837035, 
    1837036, 
    1840378, 
    1840379, 
    1843724, 
    1843725, 
    1847074, 
    1847075, 
    1850427, 
    1850428, 
    1853784, 
    1853785, 
    1857145, 
    1857146, 
    1860509, 
    1860510, 
    1863876, 
    1863877, 
    1867247, 
    1867248, 
    1870622, 
    1870623, 
    1874000, 
    1874001, 
    1877381, 
    1877382, 
    1880766, 
    1880767, 
    1884154, 
    1884155, 
    1887546, 
    1887547, 
    1890942, 
    1890943, 
    1894341, 
    1894342, 
    1897743, 
    1897744, 
    1901149, 
    1901150, 
    1904559, 
    1904560, 
    1907972, 
    1907973, 
    1911388, 
    1911389, 
    1914808, 
    1914809, 
    1918231, 
    1918232, 
    1921658, 
    1921659, 
    1925089, 
    1925090, 
    1928523, 
    1928524, 
    1931960, 
    1931961, 
    1935401, 
    1935402, 
    1938846, 
    1938847, 
    1942294, 
    1942295, 
    1945745, 
    1945746, 
    1949200, 
    1949201, 
    1952658, 
    1952659, 
    1956120, 
    1956121, 
    1959586, 
    1959587, 
    1963055, 
    1963056, 
    1966527, 
    1966528, 
    1970003, 
    1970004, 
    1973483, 
    1973484, 
    1976966, 
    1976967, 
    1980452, 
    1980453, 
    1983942, 
    1983943, 
    1987435, 
    1987436, 
    1990932, 
    1990933, 
    1994433, 
    1994434, 
    1997937, 
    1997938, 
    2001444, 
    2001445, 
    2004952, 
    2004953, 
    2008462, 
    2008463, 
    2011973, 
    2011974, 
    2015485, 
    2015486, 
    2018999, 
    2019000, 
    2022513, 
    2022514, 
    2026029, 
    2026030, 
    2029547, 
    2029548, 
    2033066, 
    2033067, 
    2036586, 
    2036587, 
    2040107, 
    2040108, 
    2043630, 
    2043631, 
    2047154, 
    2047155, 
    2050679, 
    2050680, 
    2054206, 
    2054207, 
    2057733, 
    2057734, 
    2061262, 
    2061263, 
    2064793, 
    2064794, 
    2068325, 
    2068326, 
    2071858, 
    2071859, 
    2075392, 
    2075393, 
    2078928, 
    2078929, 
    2082465, 
    2082466, 
    2086003, 
    2086004, 
    2089543, 
    2089544, 
    2093083, 
    2093084, 
    2096625, 
    2096626, 
    2100169, 
    2100170, 
    2103714, 
    2103715, 
    2107260, 
    2107261, 
    2110807, 
    2110808, 
    2114356, 
    2114357, 
    2117906, 
    2117907, 
    2121457, 
    2121458, 
    2125010, 
    2125011, 
    2128563, 
    2128564, 
    2132118, 
    2132119, 
    2135675, 
    2135676, 
    2139233, 
    2139234, 
    2142792, 
    2142793, 
    2146352, 
    2146353, 
    2149914, 
    2149915, 
    2153477, 
    2153478, 
    2157041, 
    2157042, 
    2160607, 
    2160608, 
    2164173, 
    2164174, 
    2167741, 
    2167742, 
    2171311, 
    2171312, 
    2174882, 
    2174883, 
    2178454, 
    2178455, 
    2182027, 
    2182028, 
    2185602, 
    2185603, 
    2189178, 
    2189179, 
    2192755, 
    2192756, 
    2196334, 
    2196335, 
    2199913, 
    2199914, 
    2203494, 
    2203495, 
    2207077, 
    2207078, 
    2210661, 
    2210662, 
    2214246, 
    2214247, 
    2217832, 
    2217833, 
    2221420, 
    2221421, 
    2225009, 
    2225010, 
    2228599, 
    2228600, 
    2232191, 
    2232192, 
    2235783, 
    2235784, 
    2239377, 
    2239378, 
    2242973, 
    2242974, 
    2246570, 
    2246571, 
    2250168, 
    2250169, 
    2253767, 
    2253768, 
    2257368, 
    2257369, 
    2260970, 
    2260971, 
    2264573, 
    2264574, 
    2268178, 
    2268179, 
    2271783, 
    2271784, 
    2275390, 
    2275391, 
    2278999, 
    2279000, 
    2282609, 
    2282610, 
    2286220, 
    2286221, 
    2289832, 
    2289833, 
    2293446, 
    2293447, 
    2297061, 
    2297062, 
    2300677, 
    2300678, 
    2304295, 
    2304296, 
    2307913, 
    2307914, 
    2311533, 
    2311534, 
    2315155, 
    2315156, 
    2318778, 
    2318779, 
    2322402, 
    2322403, 
    2326027, 
    2326028, 
    2329654, 
    2329655, 
    2333282, 
    2333283, 
    2336911, 
    2336912, 
    2340542, 
    2340543, 
    2344173, 
    2344174, 
    2347806, 
    2347807, 
    2351441, 
    2351442, 
    2355077, 
    2355078, 
    2358714, 
    2358715, 
    2362352, 
    2362353, 
    2365992, 
    2365993, 
    2369633, 
    2369634, 
    2373275, 
    2373276, 
    2376919, 
    2376920, 
    2380563, 
    2380564, 
    2384209, 
    2384210, 
    2387857, 
    2387858, 
    2391506, 
    2391507, 
    2395156, 
    2395157, 
    2398807, 
    2398808, 
    2402460, 
    2402461, 
    2406114, 
    2406115, 
    2409769, 
    2409770, 
    2413426, 
    2413427, 
    2417083, 
    2417084, 
    2420742, 
    2420743, 
    2424403, 
    2424404, 
    2428065, 
    2428066, 
    2431728, 
    2431729, 
    2435392, 
    2435393, 
    2439058, 
    2439059, 
    2442725, 
    2442726, 
    2446393, 
    2446394, 
    2450063, 
    2450064, 
    2453733, 
    2453734, 
    2457405, 
    2457406, 
    2461079, 
    2461080, 
    2464754, 
    2464755, 
    2468430, 
    2468431, 
    2472107, 
    2472108, 
    2475786, 
    2475787, 
    2479466, 
    2479467, 
    2483147, 
    2483148, 
    2486830, 
    2486831, 
    2490513, 
    2490514, 
    2494198, 
    2494199, 
    2497885, 
    2497886, 
    2501573, 
    2501574, 
    2505262, 
    2505263, 
    2508952, 
    2508953, 
    2512644, 
    2512645, 
    2516337, 
    2516338, 
    2520031, 
    2520032, 
    2523727, 
    2523728, 
    2527423, 
    2527424, 
    2531121, 
    2531122, 
    2534821, 
    2534822, 
    2538521, 
    2538522, 
    2542222, 
    2542223, 
    2545920, 
    2545921, 
    2549615, 
    2549616, 
    2553306, 
    2553307, 
    2556994, 
    2556995, 
    2560679, 
    2560680, 
    2564360, 
    2564361, 
    2568038, 
    2568039, 
    2571713, 
    2571714, 
    2575384, 
    2575385, 
    2579052, 
    2579053, 
    2582717, 
    2582718, 
    2586380, 
    2586381, 
    2590038, 
    2590039, 
    2593694, 
    2593695, 
    2597347, 
    2597348, 
    2600996, 
    2600997, 
    2604642, 
    2604643, 
    2608285, 
    2608286, 
    2611924, 
    2611925, 
    2615560, 
    2615561, 
    2619193, 
    2619194, 
    2622823, 
    2622824, 
    2626449, 
    2626450, 
    2630072, 
    2630073, 
    2633692, 
    2633693, 
    2637308, 
    2637309, 
    2640921, 
    2640922, 
    2644531, 
    2644532, 
    2648137, 
    2648138, 
    2651740, 
    2651741, 
    2655340, 
    2655341, 
    2658937, 
    2658938, 
    2662530, 
    2662531, 
    2666120, 
    2666121, 
    2669707, 
    2669708, 
    2673291, 
    2673292, 
    2676872, 
    2676873, 
    2680450, 
    2680451, 
    2684024, 
    2684025, 
    2687595, 
    2687596, 
    2691163, 
    2691164, 
    2694728, 
    2694729, 
    2698289, 
    2698290, 
    2701847, 
    2701848, 
    2705402, 
    2705403, 
    2708953, 
    2708954, 
    2712501, 
    2712502, 
    2716046, 
    2716047, 
    2719587, 
    2719588, 
    2723125, 
    2723126, 
    2726660, 
    2726661, 
    2730192, 
    2730193, 
    2733720, 
    2733721, 
    2737245, 
    2737246, 
    2740767, 
    2740768, 
    2744285, 
    2744286, 
    2747801, 
    2747802, 
    2751314, 
    2751315, 
    2754823, 
    2754824, 
    2758329, 
    2758330, 
    2761832, 
    2761833, 
    2765332, 
    2765333, 
    2768828, 
    2768829, 
    2772321, 
    2772322, 
    2775811, 
    2775812, 
    2779297, 
    2779298, 
    2782780, 
    2782781, 
    2786260, 
    2786261, 
    2789736, 
    2789737, 
    2793209, 
    2793210, 
    2796679, 
    2796680, 
    2800146, 
    2800147, 
    2803609, 
    2803610, 
    2807071, 
    2807072, 
    2810532, 
    2810533, 
    2813991, 
    2813992, 
    2817449, 
    2817450, 
    2820907, 
    2820908, 
    2824363, 
    2824364, 
    2827818, 
    2827819, 
    2831272, 
    2831273, 
    2834725, 
    2834726, 
    2838176, 
    2838177, 
    2841626, 
    2841627, 
    2845075, 
    2845076, 
    2848523, 
    2848524, 
    2851970, 
    2851971, 
    2855416, 
    2855417, 
    2858860, 
    2858861, 
    2862303, 
    2862304, 
    2865745, 
    2865746, 
    2869186, 
    2869187, 
    2872625, 
    2872626, 
    2876064, 
    2876065, 
    2879502, 
    2879503, 
    2882938, 
    2882939, 
    2886373, 
    2886374, 
    2889807, 
    2889808, 
    2893239, 
    2893240, 
    2896670, 
    2896671, 
    2900100, 
    2900101, 
    2903530, 
    2903531, 
    2906958, 
    2906959, 
    2910385, 
    2910386, 
    2913811, 
    2913812, 
    2917235, 
    2917236, 
    2920658, 
    2920659, 
    2924080, 
    2924081, 
    2927500, 
    2927501, 
    2930920, 
    2930921, 
    2934339, 
    2934340, 
    2937757, 
    2937758, 
    2941173, 
    2941174, 
    2944588, 
    2944589, 
    2948002, 
    2948003, 
    2951414, 
    2951415, 
    2954825, 
    2954826, 
    2958236, 
    2958237, 
    2961645, 
    2961646, 
    2965053, 
    2965054, 
    2968460, 
    2968461, 
    2971866, 
    2971867, 
    2975270, 
    2975271, 
    2978673, 
    2978674, 
    2982075, 
    2982076, 
    2985476, 
    2985477, 
    2988874, 
    2988875, 
    2992268, 
    2992269, 
    2995658, 
    2995659, 
    2999044, 
    2999045, 
    3002426, 
    3002427, 
    3005804, 
    3005805, 
    3009177, 
    3009178, 
    3012547, 
    3012548, 
    3015913, 
    3015914, 
    3019274, 
    3019275, 
    3022631, 
    3022632, 
    3025984, 
    3025985, 
    3029333, 
    3029334, 
    3032678, 
    3032679, 
    3036019, 
    3036020, 
    3039356, 
    3039357, 
    3042688, 
    3042689, 
    3046016, 
    3046017, 
    3049339, 
    3049340, 
    3052657, 
    3052658, 
    3055970, 
    3055971, 
    3059278, 
    3059279, 
    3062581, 
    3062582, 
    3065879, 
    3065880, 
    3069172, 
    3069173, 
    3072461, 
    3072462, 
    3075744, 
    3075745, 
    3079022, 
    3079023, 
    3082296, 
    3082297, 
    3085564, 
    3085565, 
    3088827, 
    3088828, 
    3092086, 
    3092087, 
    3095339, 
    3095340, 
    3098587, 
    3098588, 
    3101831, 
    3101832, 
    3105070, 
    3105071, 
    3108303, 
    3108304, 
    3111533, 
    3111534, 
    3114761, 
    3114762, 
    3117986, 
    3117987, 
    3121208, 
    3121209, 
    3124428, 
    3124429, 
    3127644, 
    3127645, 
    3130858, 
    3130859, 
    3134070, 
    3134071, 
    3137279, 
    3137280, 
    3140485, 
    3140486, 
    3143688, 
    3143689, 
    3146889, 
    3146890, 
    3150087, 
    3150088, 
    3153282, 
    3153283, 
    3156475, 
    3156476, 
    3159664, 
    3159665, 
    3162851, 
    3162852, 
    3166036, 
    3166037, 
    3169218, 
    3169219, 
    3172397, 
    3172398, 
    3175571, 
    3175572, 
    3178741, 
    3178742, 
    3181906, 
    3181907, 
    3185065, 
    3185066, 
    3188220, 
    3188221, 
    3191369, 
    3191370, 
    3194514, 
    3194515, 
    3197654, 
    3197655, 
    3200789, 
    3200790, 
    3203919, 
    3203920, 
    3207045, 
    3207046, 
    3210165, 
    3210166, 
    3213280, 
    3213281, 
    3216390, 
    3216391, 
    3219493, 
    3219494, 
    3222590, 
    3222591, 
    3225680, 
    3225681, 
    3228764, 
    3228765, 
    3231842, 
    3231843, 
    3234914, 
    3234915, 
    3237979, 
    3237980, 
    3241037, 
    3241038, 
    3244090, 
    3244091, 
    3247136, 
    3247137, 
    3250176, 
    3250177, 
    3253209, 
    3253210, 
    3256236, 
    3256237, 
    3259257, 
    3259258, 
    3262272, 
    3262273, 
    3265280, 
    3265281, 
    3268281, 
    3268282, 
    3271277, 
    3271278, 
    3274266, 
    3274267, 
    3277249, 
    3277250, 
    3280225, 
    3280226, 
    3283195, 
    3283196, 
    3286159, 
    3286160, 
    3289117, 
    3289118, 
    3292068, 
    3292069, 
    3295012, 
    3295013, 
    3297951, 
    3297952, 
    3300883, 
    3300884, 
    3303809, 
    3303810, 
    3306727, 
    3306728, 
    3309638, 
    3309639, 
    3312540, 
    3312541, 
    3315435, 
    3315436, 
    3318322, 
    3318323, 
    3321200, 
    3321201, 
    3324071, 
    3324072, 
    3326933, 
    3326934, 
    3329788, 
    3329789, 
    3332634, 
    3332635, 
    3335473, 
    3335474, 
    3338304, 
    3338305, 
    3341127, 
    3341128, 
    3343942, 
    3343943, 
    3346749, 
    3346750, 
    3349548, 
    3349549, 
    3352339, 
    3352340, 
    3355122, 
    3355123, 
    3357897, 
    3357898, 
    3360664, 
    3360665, 
    3363423, 
    3363424, 
    3366174, 
    3366175, 
    3368917, 
    3368918, 
    3371653, 
    3371654, 
    3374380, 
    3374381, 
    3377099, 
    3377100, 
    3379810, 
    3379811, 
    3382513, 
    3382514, 
    3385208, 
    3385209, 
    3387895, 
    3387896, 
    3390575, 
    3390576, 
    3393246, 
    3393247, 
    3395910, 
    3395911, 
    3398565, 
    3398566, 
    3401212, 
    3401213, 
    3403852, 
    3403853, 
    3406483, 
    3406484, 
    3409107, 
    3409108, 
    3411722, 
    3411723, 
    3414330, 
    3414331, 
    3416929, 
    3416930, 
    3419521, 
    3419522, 
    3422104, 
    3422105, 
    3424679, 
    3424680, 
    3427247, 
    3427248, 
    3429806, 
    3429807, 
    3432358, 
    3432359, 
    3434901, 
    3434902, 
    3437437, 
    3437438, 
    3439965, 
    3439966, 
    3442485, 
    3442486, 
    3444997, 
    3444998, 
    3447500, 
    3447501, 
    3449996, 
    3449997, 
    3452483, 
    3452484, 
    3454963, 
    3454964, 
    3457435, 
    3457436, 
    3459899, 
    3459900, 
    3462355, 
    3462356, 
    3464803, 
    3464804, 
    3467243, 
    3467244, 
    3469674, 
    3469675, 
    3472098, 
    3472099, 
    3474514, 
    3474515, 
    3476922, 
    3476923, 
    3479322, 
    3479323, 
    3481714, 
    3481715, 
    3484098, 
    3484099, 
    3486474, 
    3486475, 
    3488842, 
    3488843, 
    3491202, 
    3491203, 
    3493554, 
    3493555, 
    3495898, 
    3495899, 
    3498234, 
    3498235, 
    3500562, 
    3500563, 
    3502883, 
    3502884, 
    3505195, 
    3505196, 
    3507500, 
    3507501, 
    3509796, 
    3509797, 
    3512084, 
    3512085, 
    3514364, 
    3514365, 
    3516636, 
    3516637, 
    3518900, 
    3518901, 
    3521156, 
    3521157, 
    3523405, 
    3523406, 
    3525645, 
    3525646, 
    3527878, 
    3527879, 
    3530102, 
    3530103, 
    3532318, 
    3532319, 
    3534527, 
    3534528, 
    3536727, 
    3536728, 
    3538920, 
    3538921, 
    3541104, 
    3541105, 
    3543281, 
    3543282, 
    3545449, 
    3545450, 
    3547610, 
    3547611, 
    3549763, 
    3549764, 
    3551907, 
    3551908, 
    3554044, 
    3554045, 
    3556172, 
    3556173, 
    3558293, 
    3558294, 
    3560405, 
    3560406, 
    3562510, 
    3562511, 
    3564607, 
    3564608, 
    3566696, 
    3566697, 
    3568777, 
    3568778, 
    3570850, 
    3570851, 
    3572915, 
    3572916, 
    3574971, 
    3574972, 
    3577020, 
    3577021, 
    3579061, 
    3579062, 
    3581094, 
    3581095, 
    3583119, 
    3583120, 
    3585136, 
    3585137, 
    3587145, 
    3587146, 
    3589147, 
    3589148, 
    3591140, 
    3591141, 
    3593125, 
    3593126, 
    3595102, 
    3595103, 
    3597071, 
    3597072, 
    3599032, 
    3599033, 
    3600985, 
    3600986, 
    3602931, 
    3602932, 
    3604868, 
    3604869, 
    3606798, 
    3606799, 
    3608719, 
    3608720, 
    3610632, 
    3610633, 
    3612537, 
    3612538, 
    3614434, 
    3614435, 
    3616324, 
    3616325, 
    3618205, 
    3618206, 
    3620079, 
    3620080, 
    3621944, 
    3621945, 
    3623802, 
    3623803, 
    3625651, 
    3625652, 
    3627492, 
    3627493, 
    3629326, 
    3629327, 
    3631151, 
    3631152, 
    3632969, 
    3632970, 
    3634778, 
    3634779, 
    3636580, 
    3636581, 
    3638373, 
    3638374, 
    3640159, 
    3640160, 
    3641937, 
    3641938, 
    3643706, 
    3643707, 
    3645468, 
    3645469, 
    3647221, 
    3647222, 
    3648967, 
    3648968, 
    3650704, 
    3650705, 
    3652434, 
    3652435, 
    3654156, 
    3654157, 
    3655870, 
    3655871, 
    3657576, 
    3657577, 
    3659273, 
    3659274, 
    3660963, 
    3660964, 
    3662645, 
    3662646, 
    3664319, 
    3664320, 
    3665985, 
    3665986, 
    3667643, 
    3667644, 
    3669293, 
    3669294, 
    3670935, 
    3670936, 
    3672569, 
    3672570, 
    3674195, 
    3674196, 
    3675813, 
    3675814, 
    3677423, 
    3677424, 
    3679025, 
    3679026, 
    3680619, 
    3680620, 
    3682205, 
    3682206, 
    3683783, 
    3683784, 
    3685354, 
    3685355, 
    3686916, 
    3686917, 
    3688470, 
    3688471, 
    3690016, 
    3690017, 
    3691554, 
    3691555, 
    3693084, 
    3693085, 
    3694606, 
    3694607, 
    3696121, 
    3696122, 
    3697627, 
    3697628, 
    3699126, 
    3699127, 
    3700616, 
    3700617, 
    3702098, 
    3702099, 
    3703572, 
    3703573, 
    3705038, 
    3705039, 
    3706497, 
    3706498, 
    3707947, 
    3707948, 
    3709390, 
    3709391, 
    3710824, 
    3710825, 
    3712251, 
    3712252, 
    3713669, 
    3713670, 
    3715079, 
    3715080, 
    3716482, 
    3716483, 
    3717876, 
    3717877, 
    3719263, 
    3719264, 
    3720641, 
    3720642, 
    3722012, 
    3722013, 
    3723375, 
    3723376, 
    3724730, 
    3724731, 
    3726077, 
    3726078, 
    3727416, 
    3727417, 
    3728747, 
    3728748, 
    3730069, 
    3730070, 
    3731384, 
    3731385, 
    3732691, 
    3732692, 
    3733990, 
    3733991, 
    3735281, 
    3735282, 
    3736564, 
    3736565, 
    3737839, 
    3737840, 
    3739106, 
    3739107, 
    3740365, 
    3740366, 
    3741616, 
    3741617, 
    3742859, 
    3742860, 
    3744094, 
    3744095, 
    3745321, 
    3745322, 
    3746540, 
    3746541, 
    3747751, 
    3747752, 
    3748954, 
    3748955, 
    3750150, 
    3750151, 
    3751337, 
    3751338, 
    3752516, 
    3752517, 
    3753687, 
    3753688, 
    3754850, 
    3754851, 
    3756005, 
    3756006, 
    3757152, 
    3757153, 
    3758292, 
    3758293, 
    3759423, 
    3759424, 
    3760547, 
    3760548, 
    3761662, 
    3761663, 
    3762769, 
    3762770, 
    3763868, 
    3763869, 
    3764959, 
    3764960, 
    3766043, 
    3766044, 
    3767118, 
    3767119, 
    3768186, 
    3768187, 
    3769245, 
    3769246, 
    3770297, 
    3770298, 
    3771341, 
    3771342, 
    3772376, 
    3772377, 
    3773404, 
    3773405, 
    3774423, 
    3774424, 
    3775435, 
    3775436, 
    3776438, 
    3776439, 
    3777434, 
    3777435, 
    3778422, 
    3778423, 
    3779394, 
    3779395, 
    3780318, 
    3780319, 
    3781191, 
    3781192, 
    3782017, 
    3782018, 
    3782793, 
    3782794, 
    3783521, 
    3783522, 
    3784198, 
    3784199, 
    3784828, 
    3784829, 
    3785408, 
    3785409, 
    3785939, 
    3785940, 
    3786420, 
    3786421, 
    3786853, 
    3786854, 
    3787237, 
    3787238, 
    3787571, 
    3787572, 
    3787857, 
    3787858, 
    3788094, 
    3788095, 
    3788282, 
    3788283, 
    3788420, 
    3788421, 
    3788510, 
    3788511 ;

 runlens = 
    1, 
    1, 
    2, 
    1, 
    5, 
    1, 
    7, 
    1, 
    9, 
    1, 
    11, 
    1, 
    14, 
    1, 
    16, 
    1, 
    18, 
    1, 
    20, 
    1, 
    23, 
    1, 
    26, 
    1, 
    28, 
    1, 
    30, 
    1, 
    33, 
    1, 
    35, 
    1, 
    37, 
    1, 
    39, 
    1, 
    42, 
    1, 
    44, 
    1, 
    46, 
    1, 
    48, 
    1, 
    51, 
    1, 
    53, 
    1, 
    55, 
    1, 
    58, 
    1, 
    60, 
    1, 
    62, 
    1, 
    64, 
    1, 
    67, 
    1, 
    69, 
    1, 
    71, 
    1, 
    73, 
    1, 
    76, 
    1, 
    78, 
    1, 
    80, 
    1, 
    82, 
    1, 
    85, 
    1, 
    87, 
    1, 
    89, 
    1, 
    91, 
    1, 
    95, 
    1, 
    97, 
    1, 
    99, 
    1, 
    101, 
    1, 
    104, 
    1, 
    106, 
    1, 
    108, 
    1, 
    110, 
    1, 
    113, 
    1, 
    115, 
    1, 
    117, 
    1, 
    120, 
    1, 
    122, 
    1, 
    124, 
    1, 
    126, 
    1, 
    129, 
    1, 
    131, 
    1, 
    133, 
    1, 
    135, 
    1, 
    138, 
    1, 
    140, 
    1, 
    142, 
    1, 
    144, 
    1, 
    147, 
    1, 
    149, 
    1, 
    151, 
    1, 
    153, 
    1, 
    156, 
    1, 
    158, 
    1, 
    160, 
    1, 
    163, 
    1, 
    166, 
    1, 
    168, 
    1, 
    170, 
    1, 
    173, 
    1, 
    175, 
    1, 
    177, 
    1, 
    179, 
    1, 
    182, 
    1, 
    184, 
    1, 
    186, 
    1, 
    188, 
    1, 
    191, 
    1, 
    193, 
    1, 
    195, 
    1, 
    197, 
    1, 
    200, 
    1, 
    202, 
    1, 
    204, 
    1, 
    206, 
    1, 
    209, 
    1, 
    211, 
    1, 
    213, 
    1, 
    215, 
    1, 
    218, 
    1, 
    220, 
    1, 
    222, 
    1, 
    224, 
    1, 
    227, 
    1, 
    229, 
    1, 
    231, 
    1, 
    235, 
    1, 
    237, 
    1, 
    239, 
    1, 
    241, 
    1, 
    244, 
    1, 
    246, 
    1, 
    248, 
    1, 
    250, 
    1, 
    253, 
    1, 
    255, 
    1, 
    257, 
    1, 
    259, 
    1, 
    262, 
    1, 
    264, 
    1, 
    266, 
    1, 
    268, 
    1, 
    271, 
    1, 
    273, 
    1, 
    275, 
    1, 
    277, 
    1, 
    280, 
    1, 
    282, 
    1, 
    284, 
    1, 
    287, 
    1, 
    289, 
    1, 
    291, 
    1, 
    293, 
    1, 
    296, 
    1, 
    298, 
    1, 
    300, 
    1, 
    303, 
    1, 
    306, 
    1, 
    308, 
    1, 
    310, 
    1, 
    312, 
    1, 
    315, 
    1, 
    317, 
    1, 
    319, 
    1, 
    321, 
    1, 
    324, 
    1, 
    326, 
    1, 
    328, 
    1, 
    330, 
    1, 
    333, 
    1, 
    335, 
    1, 
    337, 
    1, 
    339, 
    1, 
    342, 
    1, 
    344, 
    1, 
    346, 
    1, 
    349, 
    1, 
    351, 
    1, 
    353, 
    1, 
    355, 
    1, 
    358, 
    1, 
    360, 
    1, 
    362, 
    1, 
    364, 
    1, 
    367, 
    1, 
    369, 
    1, 
    371, 
    1, 
    374, 
    1, 
    377, 
    1, 
    379, 
    1, 
    381, 
    1, 
    383, 
    1, 
    386, 
    1, 
    388, 
    1, 
    390, 
    1, 
    392, 
    1, 
    395, 
    1, 
    397, 
    1, 
    399, 
    1, 
    402, 
    1, 
    404, 
    1, 
    406, 
    1, 
    408, 
    1, 
    411, 
    1, 
    413, 
    1, 
    415, 
    1, 
    417, 
    1, 
    420, 
    1, 
    422, 
    1, 
    424, 
    1, 
    426, 
    1, 
    429, 
    1, 
    431, 
    1, 
    433, 
    1, 
    435, 
    1, 
    438, 
    1, 
    440, 
    1, 
    443, 
    1, 
    445, 
    1, 
    448, 
    1, 
    450, 
    1, 
    452, 
    1, 
    454, 
    1, 
    457, 
    1, 
    459, 
    1, 
    461, 
    1, 
    464, 
    1, 
    466, 
    1, 
    468, 
    1, 
    470, 
    1, 
    473, 
    1, 
    475, 
    1, 
    477, 
    1, 
    479, 
    1, 
    482, 
    1, 
    484, 
    1, 
    486, 
    1, 
    488, 
    1, 
    491, 
    1, 
    493, 
    1, 
    495, 
    1, 
    497, 
    1, 
    500, 
    1, 
    502, 
    1, 
    504, 
    1, 
    506, 
    1, 
    509, 
    1, 
    512, 
    1, 
    514, 
    1, 
    517, 
    1, 
    519, 
    1, 
    521, 
    1, 
    523, 
    1, 
    526, 
    1, 
    528, 
    1, 
    530, 
    1, 
    532, 
    1, 
    535, 
    1, 
    537, 
    1, 
    539, 
    1, 
    541, 
    1, 
    544, 
    1, 
    546, 
    1, 
    548, 
    1, 
    550, 
    1, 
    553, 
    1, 
    555, 
    1, 
    557, 
    1, 
    559, 
    1, 
    562, 
    1, 
    564, 
    1, 
    566, 
    1, 
    568, 
    1, 
    571, 
    1, 
    573, 
    1, 
    575, 
    1, 
    578, 
    1, 
    581, 
    1, 
    583, 
    1, 
    585, 
    1, 
    588, 
    1, 
    590, 
    1, 
    592, 
    1, 
    594, 
    1, 
    597, 
    1, 
    599, 
    1, 
    601, 
    1, 
    603, 
    1, 
    606, 
    1, 
    608, 
    1, 
    610, 
    1, 
    612, 
    1, 
    615, 
    1, 
    617, 
    1, 
    619, 
    1, 
    621, 
    1, 
    624, 
    1, 
    626, 
    1, 
    628, 
    1, 
    631, 
    1, 
    633, 
    1, 
    635, 
    1, 
    637, 
    1, 
    640, 
    1, 
    642, 
    1, 
    644, 
    1, 
    646, 
    1, 
    649, 
    1, 
    652, 
    1, 
    654, 
    1, 
    656, 
    1, 
    659, 
    1, 
    661, 
    1, 
    663, 
    1, 
    665, 
    1, 
    668, 
    1, 
    670, 
    1, 
    672, 
    1, 
    674, 
    1, 
    677, 
    1, 
    679, 
    1, 
    681, 
    1, 
    683, 
    1, 
    686, 
    1, 
    688, 
    1, 
    690, 
    1, 
    693, 
    1, 
    695, 
    1, 
    697, 
    1, 
    699, 
    1, 
    702, 
    1, 
    704, 
    1, 
    706, 
    1, 
    708, 
    1, 
    711, 
    1, 
    713, 
    1, 
    715, 
    1, 
    717, 
    1, 
    720, 
    1, 
    723, 
    1, 
    725, 
    1, 
    727, 
    1, 
    730, 
    1, 
    732, 
    1, 
    734, 
    1, 
    736, 
    1, 
    739, 
    1, 
    741, 
    1, 
    743, 
    1, 
    746, 
    1, 
    748, 
    1, 
    750, 
    1, 
    752, 
    1, 
    755, 
    1, 
    757, 
    1, 
    759, 
    1, 
    761, 
    1, 
    764, 
    1, 
    766, 
    1, 
    768, 
    1, 
    770, 
    1, 
    773, 
    1, 
    775, 
    1, 
    777, 
    1, 
    779, 
    1, 
    782, 
    1, 
    784, 
    1, 
    786, 
    1, 
    788, 
    1, 
    792, 
    1, 
    794, 
    1, 
    796, 
    1, 
    798, 
    1, 
    801, 
    1, 
    803, 
    1, 
    805, 
    1, 
    808, 
    1, 
    810, 
    1, 
    812, 
    1, 
    814, 
    1, 
    817, 
    1, 
    819, 
    1, 
    821, 
    1, 
    823, 
    1, 
    826, 
    1, 
    828, 
    1, 
    830, 
    1, 
    832, 
    1, 
    835, 
    1, 
    837, 
    1, 
    839, 
    1, 
    841, 
    1, 
    844, 
    1, 
    846, 
    1, 
    848, 
    1, 
    850, 
    1, 
    853, 
    1, 
    855, 
    1, 
    857, 
    1, 
    861, 
    1, 
    863, 
    1, 
    865, 
    1, 
    867, 
    1, 
    870, 
    1, 
    872, 
    1, 
    874, 
    1, 
    876, 
    1, 
    879, 
    1, 
    881, 
    1, 
    883, 
    1, 
    885, 
    1, 
    888, 
    1, 
    890, 
    1, 
    892, 
    1, 
    894, 
    1, 
    897, 
    1, 
    899, 
    1, 
    901, 
    1, 
    903, 
    1, 
    906, 
    1, 
    908, 
    1, 
    910, 
    1, 
    912, 
    1, 
    915, 
    1, 
    917, 
    1, 
    919, 
    1, 
    921, 
    1, 
    924, 
    1, 
    926, 
    1, 
    928, 
    1, 
    932, 
    1, 
    934, 
    1, 
    936, 
    1, 
    938, 
    1, 
    941, 
    1, 
    943, 
    1, 
    945, 
    1, 
    947, 
    1, 
    950, 
    1, 
    952, 
    1, 
    954, 
    1, 
    956, 
    1, 
    959, 
    1, 
    961, 
    1, 
    963, 
    1, 
    965, 
    1, 
    968, 
    1, 
    970, 
    1, 
    972, 
    1, 
    975, 
    1, 
    977, 
    1, 
    979, 
    1, 
    981, 
    1, 
    984, 
    1, 
    986, 
    1, 
    988, 
    1, 
    990, 
    1, 
    993, 
    1, 
    995, 
    1, 
    997, 
    1, 
    1000, 
    1, 
    1003, 
    1, 
    1005, 
    1, 
    1007, 
    1, 
    1009, 
    1, 
    1012, 
    1, 
    1014, 
    1, 
    1016, 
    1, 
    1018, 
    1, 
    1021, 
    1, 
    1023, 
    1, 
    1025, 
    1, 
    1027, 
    1, 
    1030, 
    1, 
    1032, 
    1, 
    1034, 
    1, 
    1036, 
    1, 
    1039, 
    1, 
    1041, 
    1, 
    1043, 
    1, 
    1046, 
    1, 
    1048, 
    1, 
    1050, 
    1, 
    1052, 
    1, 
    1055, 
    1, 
    1057, 
    1, 
    1059, 
    1, 
    1061, 
    1, 
    1064, 
    1, 
    1066, 
    1, 
    1068, 
    1, 
    1071, 
    1, 
    1074, 
    1, 
    1076, 
    1, 
    1078, 
    1, 
    1080, 
    1, 
    1083, 
    1, 
    1085, 
    1, 
    1087, 
    1, 
    1090, 
    1, 
    1092, 
    1, 
    1094, 
    1, 
    1096, 
    1, 
    1099, 
    1, 
    1101, 
    1, 
    1103, 
    1, 
    1105, 
    1, 
    1108, 
    1, 
    1110, 
    1, 
    1112, 
    1, 
    1114, 
    1, 
    1117, 
    1, 
    1119, 
    1, 
    1121, 
    1, 
    1123, 
    1, 
    1126, 
    1, 
    1128, 
    1, 
    1130, 
    1, 
    1132, 
    1, 
    1135, 
    1, 
    1137, 
    1, 
    1140, 
    1, 
    1142, 
    1, 
    1145, 
    1, 
    1147, 
    1, 
    1149, 
    1, 
    1152, 
    1, 
    1154, 
    1, 
    1156, 
    1, 
    1158, 
    1, 
    1161, 
    1, 
    1163, 
    1, 
    1165, 
    1, 
    1167, 
    1, 
    1170, 
    1, 
    1172, 
    1, 
    1174, 
    1, 
    1176, 
    1, 
    1179, 
    1, 
    1181, 
    1, 
    1183, 
    1, 
    1185, 
    1, 
    1188, 
    1, 
    1190, 
    1, 
    1192, 
    1, 
    1194, 
    1, 
    1197, 
    1, 
    1199, 
    1, 
    1201, 
    1, 
    1204, 
    1, 
    1206, 
    1, 
    1209, 
    1, 
    1211, 
    1, 
    1214, 
    1, 
    1216, 
    1, 
    1218, 
    1, 
    1220, 
    1, 
    1223, 
    1, 
    1225, 
    1, 
    1227, 
    1, 
    1229, 
    1, 
    1232, 
    1, 
    1234, 
    1, 
    1236, 
    1, 
    1238, 
    1, 
    1241, 
    1, 
    1243, 
    1, 
    1245, 
    1, 
    1247, 
    1, 
    1250, 
    1, 
    1252, 
    1, 
    1254, 
    1, 
    1256, 
    1, 
    1259, 
    1, 
    1261, 
    1, 
    1263, 
    1, 
    1266, 
    1, 
    1268, 
    1, 
    1270, 
    1, 
    1272, 
    1, 
    1275, 
    1, 
    1277, 
    1, 
    1280, 
    1, 
    1282, 
    1, 
    1285, 
    1, 
    1287, 
    1, 
    1289, 
    1, 
    1291, 
    1, 
    1294, 
    1, 
    1296, 
    1, 
    1298, 
    1, 
    1300, 
    1, 
    1303, 
    1, 
    1305, 
    1, 
    1307, 
    1, 
    1309, 
    1, 
    1312, 
    1, 
    1314, 
    1, 
    1316, 
    1, 
    1319, 
    1, 
    1321, 
    1, 
    1323, 
    1, 
    1325, 
    1, 
    1328, 
    1, 
    1330, 
    1, 
    1332, 
    1, 
    1334, 
    1, 
    1337, 
    1, 
    1339, 
    1, 
    1341, 
    1, 
    1343, 
    1, 
    1346, 
    1, 
    1349, 
    1, 
    1351, 
    1, 
    1353, 
    1, 
    1356, 
    1, 
    1358, 
    1, 
    1360, 
    1, 
    1362, 
    1, 
    1365, 
    1, 
    1367, 
    1, 
    1369, 
    1, 
    1371, 
    1, 
    1374, 
    1, 
    1376, 
    1, 
    1378, 
    1, 
    1381, 
    1, 
    1383, 
    1, 
    1385, 
    1, 
    1387, 
    1, 
    1390, 
    1, 
    1392, 
    1, 
    1394, 
    1, 
    1396, 
    1, 
    1399, 
    1, 
    1401, 
    1, 
    1403, 
    1, 
    1405, 
    1, 
    1408, 
    1, 
    1410, 
    1, 
    1412, 
    1, 
    1414, 
    1, 
    1417, 
    1, 
    1420, 
    1, 
    1422, 
    1, 
    1424, 
    1, 
    1427, 
    1, 
    1429, 
    1, 
    1431, 
    1, 
    1434, 
    1, 
    1436, 
    1, 
    1438, 
    1, 
    1440, 
    1, 
    1443, 
    1, 
    1445, 
    1, 
    1447, 
    1, 
    1449, 
    1, 
    1452, 
    1, 
    1454, 
    1, 
    1456, 
    1, 
    1458, 
    1, 
    1461, 
    1, 
    1463, 
    1, 
    1465, 
    1, 
    1467, 
    1, 
    1470, 
    1, 
    1472, 
    1, 
    1474, 
    1, 
    1476, 
    1, 
    1479, 
    1, 
    1481, 
    1, 
    1483, 
    1, 
    1485, 
    1, 
    1489, 
    1, 
    1491, 
    1, 
    1493, 
    1, 
    1496, 
    1, 
    1498, 
    1, 
    1500, 
    1, 
    1502, 
    1, 
    1505, 
    1, 
    1507, 
    1, 
    1509, 
    1, 
    1511, 
    1, 
    1514, 
    1, 
    1516, 
    1, 
    1518, 
    1, 
    1520, 
    1, 
    1523, 
    1, 
    1525, 
    1, 
    1527, 
    1, 
    1531, 
    1, 
    1536, 
    1, 
    1541, 
    1, 
    1545, 
    1, 
    1550, 
    1, 
    1554, 
    1, 
    1559, 
    1, 
    1563, 
    1, 
    1568, 
    1, 
    1573, 
    1, 
    1577, 
    1, 
    1582, 
    1, 
    1587, 
    1, 
    1592, 
    1, 
    1596, 
    1, 
    1601, 
    1, 
    1606, 
    1, 
    1610, 
    1, 
    1615, 
    1, 
    1619, 
    1, 
    1624, 
    1, 
    1628, 
    1, 
    1633, 
    1, 
    1637, 
    1, 
    1642, 
    1, 
    1647, 
    1, 
    1651, 
    1, 
    1656, 
    1, 
    1660, 
    1, 
    1665, 
    1, 
    1669, 
    1, 
    1674, 
    1, 
    1679, 
    1, 
    1683, 
    1, 
    1688, 
    1, 
    1692, 
    1, 
    1697, 
    1, 
    1701, 
    1, 
    1706, 
    1, 
    1711, 
    1, 
    1715, 
    1, 
    1720, 
    1, 
    1724, 
    1, 
    1730, 
    1, 
    1734, 
    1, 
    1739, 
    1, 
    1744, 
    1, 
    1748, 
    1, 
    1753, 
    1, 
    1757, 
    1, 
    1762, 
    1, 
    1766, 
    1, 
    1771, 
    1, 
    1775, 
    1, 
    1780, 
    1, 
    1785, 
    1, 
    1789, 
    1, 
    1794, 
    1, 
    1798, 
    1, 
    1803, 
    1, 
    1807, 
    1, 
    1812, 
    1, 
    1817, 
    1, 
    1821, 
    1, 
    1826, 
    1, 
    1830, 
    1, 
    1835, 
    1, 
    1839, 
    1, 
    1844, 
    1, 
    1849, 
    1, 
    1853, 
    1, 
    1858, 
    1, 
    1862, 
    1, 
    1868, 
    1, 
    1872, 
    1, 
    1877, 
    1, 
    1882, 
    1, 
    1886, 
    1, 
    1891, 
    1, 
    1895, 
    1, 
    1900, 
    1, 
    1904, 
    1, 
    1909, 
    1, 
    1913, 
    1, 
    1918, 
    1, 
    1922, 
    1, 
    1927, 
    1, 
    1932, 
    1, 
    1936, 
    1, 
    1941, 
    1, 
    1945, 
    1, 
    1950, 
    1, 
    1955, 
    1, 
    1959, 
    1, 
    1964, 
    1, 
    1968, 
    1, 
    1973, 
    1, 
    1977, 
    1, 
    1982, 
    1, 
    1987, 
    1, 
    1991, 
    1, 
    1996, 
    1, 
    2000, 
    1, 
    2005, 
    1, 
    2010, 
    1, 
    2015, 
    1, 
    2020, 
    1, 
    2024, 
    1, 
    2029, 
    1, 
    2033, 
    1, 
    2038, 
    1, 
    2042, 
    1, 
    2047, 
    1, 
    2051, 
    1, 
    2056, 
    1, 
    2061, 
    1, 
    2065, 
    1, 
    2070, 
    1, 
    2074, 
    1, 
    2079, 
    1, 
    2083, 
    1, 
    2088, 
    1, 
    2093, 
    1, 
    2097, 
    1, 
    2102, 
    1, 
    2106, 
    1, 
    2111, 
    1, 
    2115, 
    1, 
    2120, 
    1, 
    2125, 
    1, 
    2129, 
    1, 
    2134, 
    1, 
    2138, 
    1, 
    2143, 
    1, 
    2148, 
    1, 
    2153, 
    1, 
    2158, 
    1, 
    2162, 
    1, 
    2167, 
    1, 
    2171, 
    1, 
    2176, 
    1, 
    2180, 
    1, 
    2185, 
    1, 
    2189, 
    1, 
    2194, 
    1, 
    2199, 
    1, 
    2203, 
    1, 
    2208, 
    1, 
    2212, 
    1, 
    2217, 
    1, 
    2221, 
    1, 
    2226, 
    1, 
    2231, 
    1, 
    2235, 
    1, 
    2240, 
    1, 
    2244, 
    1, 
    2249, 
    1, 
    2253, 
    1, 
    2258, 
    1, 
    2263, 
    1, 
    2267, 
    1, 
    2272, 
    1, 
    2276, 
    1, 
    2281, 
    1, 
    2286, 
    1, 
    2291, 
    1, 
    2296, 
    1, 
    2300, 
    1, 
    2305, 
    1, 
    2309, 
    1, 
    2314, 
    1, 
    2318, 
    1, 
    2323, 
    1, 
    2327, 
    1, 
    2332, 
    1, 
    2336, 
    1, 
    2341, 
    1, 
    2346, 
    1, 
    2350, 
    1, 
    2355, 
    1, 
    2359, 
    1, 
    2364, 
    1, 
    2369, 
    1, 
    2373, 
    1, 
    2378, 
    1, 
    2382, 
    1, 
    2387, 
    1, 
    2391, 
    1, 
    2396, 
    1, 
    2401, 
    1, 
    2405, 
    1, 
    2410, 
    1, 
    2414, 
    1, 
    2419, 
    1, 
    2423, 
    1, 
    2429, 
    1, 
    2434, 
    1, 
    2438, 
    1, 
    2443, 
    1, 
    2447, 
    1, 
    2449, 
    1, 
    2451, 
    1, 
    2453, 
    1, 
    2454, 
    1, 
    2456, 
    1, 
    2458, 
    1, 
    2459, 
    1, 
    2461, 
    1, 
    2463, 
    1, 
    2465, 
    1, 
    2466, 
    1, 
    2468, 
    1, 
    2470, 
    1, 
    2471, 
    1, 
    2473, 
    1, 
    2475, 
    1, 
    2476, 
    1, 
    2478, 
    1, 
    2480, 
    1, 
    2482, 
    1, 
    2483, 
    1, 
    2485, 
    1, 
    2487, 
    1, 
    2488, 
    1, 
    2490, 
    1, 
    2493, 
    1, 
    2494, 
    1, 
    2496, 
    1, 
    2498, 
    1, 
    2500, 
    1, 
    2501, 
    1, 
    2503, 
    1, 
    2505, 
    1, 
    2506, 
    1, 
    2508, 
    1, 
    2510, 
    1, 
    2511, 
    1, 
    2513, 
    1, 
    2515, 
    1, 
    2517, 
    1, 
    2518, 
    1, 
    2520, 
    1, 
    2522, 
    1, 
    2523, 
    1, 
    2525, 
    1, 
    2527, 
    1, 
    2528, 
    1, 
    2530, 
    1, 
    2532, 
    1, 
    2534, 
    1, 
    2535, 
    1, 
    2537, 
    1, 
    2539, 
    1, 
    2540, 
    1, 
    2542, 
    1, 
    2544, 
    1, 
    2546, 
    1, 
    2548, 
    1, 
    2550, 
    1, 
    2552, 
    1, 
    2553, 
    1, 
    2555, 
    1, 
    2557, 
    1, 
    2558, 
    1, 
    2560, 
    1, 
    2562, 
    1, 
    2563, 
    1, 
    2565, 
    1, 
    2567, 
    1, 
    2569, 
    1, 
    2570, 
    1, 
    2572, 
    1, 
    2574, 
    1, 
    2575, 
    1, 
    2577, 
    1, 
    2579, 
    1, 
    2580, 
    1, 
    2582, 
    1, 
    2584, 
    1, 
    2586, 
    1, 
    2587, 
    1, 
    2589, 
    1, 
    2591, 
    1, 
    2592, 
    1, 
    2594, 
    1, 
    2596, 
    1, 
    2598, 
    1, 
    2600, 
    1, 
    2602, 
    1, 
    2604, 
    1, 
    2605, 
    1, 
    2607, 
    1, 
    2609, 
    1, 
    2610, 
    1, 
    2612, 
    1, 
    2614, 
    1, 
    2615, 
    1, 
    2617, 
    1, 
    2619, 
    1, 
    2620, 
    1, 
    2622, 
    1, 
    2624, 
    1, 
    2626, 
    1, 
    2627, 
    1, 
    2629, 
    1, 
    2631, 
    1, 
    2632, 
    1, 
    2634, 
    1, 
    2636, 
    1, 
    2637, 
    1, 
    2639, 
    1, 
    2641, 
    1, 
    2643, 
    1, 
    2644, 
    1, 
    2646, 
    1, 
    2648, 
    1, 
    2650, 
    1, 
    2652, 
    1, 
    2654, 
    1, 
    2655, 
    1, 
    2657, 
    1, 
    2659, 
    1, 
    2661, 
    1, 
    2662, 
    1, 
    2664, 
    1, 
    2666, 
    1, 
    2667, 
    1, 
    2669, 
    1, 
    2671, 
    1, 
    2672, 
    1, 
    2674, 
    1, 
    2676, 
    1, 
    2678, 
    1, 
    2679, 
    1, 
    2681, 
    1, 
    2683, 
    1, 
    2684, 
    1, 
    2686, 
    1, 
    2688, 
    1, 
    2689, 
    1, 
    2691, 
    1, 
    2693, 
    1, 
    2695, 
    1, 
    2696, 
    1, 
    2698, 
    1, 
    2700, 
    1, 
    2702, 
    1, 
    2706, 
    1, 
    2709, 
    1, 
    2712, 
    1, 
    2716, 
    1, 
    2720, 
    1, 
    2724, 
    1, 
    2726, 
    1, 
    2730, 
    1, 
    2734, 
    1, 
    2737, 
    1, 
    2741, 
    1, 
    2744, 
    1, 
    2747, 
    1, 
    2751, 
    1, 
    2755, 
    1, 
    2759, 
    1, 
    2761, 
    1, 
    2765, 
    1, 
    2769, 
    1, 
    2772, 
    1, 
    2776, 
    1, 
    2779, 
    1, 
    2782, 
    1, 
    2786, 
    1, 
    2790, 
    1, 
    2793, 
    1, 
    2796, 
    1, 
    2800, 
    1, 
    2804, 
    1, 
    2807, 
    1, 
    2810, 
    1, 
    2814, 
    1, 
    2817, 
    1, 
    2821, 
    1, 
    2825, 
    1, 
    2828, 
    1, 
    2831, 
    1, 
    2835, 
    1, 
    2839, 
    1, 
    2842, 
    1, 
    2845, 
    1, 
    2849, 
    1, 
    2852, 
    1, 
    2856, 
    1, 
    2860, 
    1, 
    2863, 
    1, 
    2866, 
    1, 
    2870, 
    1, 
    2874, 
    1, 
    2877, 
    1, 
    2880, 
    1, 
    2884, 
    1, 
    2887, 
    1, 
    2891, 
    1, 
    2895, 
    1, 
    2898, 
    1, 
    2901, 
    1, 
    2905, 
    1, 
    2909, 
    1, 
    2912, 
    1, 
    2915, 
    1, 
    2919, 
    1, 
    2922, 
    1, 
    2926, 
    1, 
    2930, 
    1, 
    2933, 
    1, 
    2936, 
    1, 
    2940, 
    1, 
    2944, 
    1, 
    2947, 
    1, 
    2950, 
    1, 
    2954, 
    1, 
    2957, 
    1, 
    2961, 
    1, 
    2965, 
    1, 
    2968, 
    1, 
    2971, 
    1, 
    2975, 
    1, 
    2979, 
    1, 
    2982, 
    1, 
    2985, 
    1, 
    2989, 
    1, 
    2992, 
    1, 
    2996, 
    1, 
    3000, 
    1, 
    3003, 
    1, 
    3006, 
    1, 
    3010, 
    1, 
    3014, 
    1, 
    3017, 
    1, 
    3020, 
    1, 
    3024, 
    1, 
    3027, 
    1, 
    3031, 
    1, 
    3034, 
    1, 
    3038, 
    1, 
    3041, 
    1, 
    3045, 
    1, 
    3049, 
    1, 
    3051, 
    1, 
    3055, 
    1, 
    3059, 
    1, 
    3062, 
    1, 
    3066, 
    1, 
    3069, 
    1, 
    3073, 
    1, 
    3076, 
    1, 
    3080, 
    1, 
    3084, 
    1, 
    3086, 
    1, 
    3090, 
    1, 
    3094, 
    1, 
    3097, 
    1, 
    3101, 
    1, 
    3104, 
    1, 
    3108, 
    1, 
    3111, 
    1, 
    3115, 
    1, 
    3119, 
    1, 
    3121, 
    1, 
    3125, 
    1, 
    3129, 
    1, 
    3132, 
    1, 
    3136, 
    1, 
    3139, 
    1, 
    3143, 
    1, 
    3146, 
    1, 
    3150, 
    1, 
    3154, 
    1, 
    3156, 
    1, 
    3160, 
    1, 
    3164, 
    1, 
    3167, 
    1, 
    3171, 
    1, 
    3174, 
    1, 
    3178, 
    1, 
    3181, 
    1, 
    3185, 
    1, 
    3189, 
    1, 
    3191, 
    1, 
    3195, 
    1, 
    3199, 
    1, 
    3202, 
    1, 
    3206, 
    1, 
    3209, 
    1, 
    3213, 
    1, 
    3216, 
    1, 
    3220, 
    1, 
    3224, 
    1, 
    3226, 
    1, 
    3230, 
    1, 
    3234, 
    1, 
    3237, 
    1, 
    3241, 
    1, 
    3244, 
    1, 
    3248, 
    1, 
    3251, 
    1, 
    3255, 
    1, 
    3259, 
    1, 
    3261, 
    1, 
    3265, 
    1, 
    3269, 
    1, 
    3272, 
    1, 
    3275, 
    1, 
    3279, 
    1, 
    3282, 
    1, 
    3286, 
    1, 
    3290, 
    1, 
    3293, 
    1, 
    3296, 
    1, 
    3300, 
    1, 
    3304, 
    1, 
    3307, 
    1, 
    3310, 
    1, 
    3314, 
    1, 
    3317, 
    1, 
    3321, 
    1, 
    3325, 
    1, 
    3328, 
    1, 
    3331, 
    1, 
    3335, 
    1, 
    3339, 
    1, 
    3342, 
    1, 
    3345, 
    1, 
    3349, 
    1, 
    3352, 
    1, 
    3356, 
    1, 
    3360, 
    1, 
    3363, 
    1, 
    3366, 
    1, 
    3370, 
    1, 
    3374, 
    1, 
    3377, 
    1, 
    3380, 
    1, 
    3384, 
    1, 
    3387, 
    1, 
    3391, 
    1, 
    3395, 
    1, 
    3398, 
    1, 
    3401, 
    1, 
    3405, 
    1, 
    3409, 
    1, 
    3412, 
    1, 
    3415, 
    1, 
    3419, 
    1, 
    3422, 
    1, 
    3426, 
    1, 
    3430, 
    1, 
    3433, 
    1, 
    3436, 
    1, 
    3440, 
    1, 
    3444, 
    1, 
    3447, 
    1, 
    3450, 
    1, 
    3454, 
    1, 
    3457, 
    1, 
    3461, 
    1, 
    3465, 
    1, 
    3468, 
    1, 
    3471, 
    1, 
    3475, 
    1, 
    3479, 
    1, 
    3482, 
    1, 
    3485, 
    1, 
    3489, 
    1, 
    3492, 
    1, 
    3496, 
    1, 
    3500, 
    1, 
    3503, 
    1, 
    3506, 
    1, 
    3507, 
    1, 
    3509, 
    1, 
    3510, 
    1, 
    3511, 
    1, 
    3513, 
    1, 
    3513, 
    1, 
    3515, 
    1, 
    3517, 
    1, 
    3518, 
    1, 
    3519, 
    1, 
    3520, 
    1, 
    3522, 
    1, 
    3523, 
    1, 
    3524, 
    1, 
    3526, 
    1, 
    3526, 
    1, 
    3528, 
    1, 
    3530, 
    1, 
    3531, 
    1, 
    3532, 
    1, 
    3533, 
    1, 
    3535, 
    1, 
    3536, 
    1, 
    3537, 
    1, 
    3539, 
    1, 
    3539, 
    1, 
    3541, 
    1, 
    3543, 
    1, 
    3544, 
    1, 
    3545, 
    1, 
    3546, 
    1, 
    3548, 
    1, 
    3549, 
    1, 
    3550, 
    1, 
    3552, 
    1, 
    3552, 
    1, 
    3554, 
    1, 
    3556, 
    1, 
    3557, 
    1, 
    3558, 
    1, 
    3559, 
    1, 
    3561, 
    1, 
    3562, 
    1, 
    3563, 
    1, 
    3565, 
    1, 
    3565, 
    1, 
    3567, 
    1, 
    3569, 
    1, 
    3570, 
    1, 
    3571, 
    1, 
    3572, 
    1, 
    3574, 
    1, 
    3575, 
    1, 
    3576, 
    1, 
    3578, 
    1, 
    3578, 
    1, 
    3580, 
    1, 
    3582, 
    1, 
    3583, 
    1, 
    3584, 
    1, 
    3585, 
    1, 
    3587, 
    1, 
    3588, 
    1, 
    3589, 
    1, 
    3591, 
    1, 
    3591, 
    1, 
    3593, 
    1, 
    3595, 
    1, 
    3596, 
    1, 
    3597, 
    1, 
    3598, 
    1, 
    3600, 
    1, 
    3601, 
    1, 
    3602, 
    1, 
    3604, 
    1, 
    3604, 
    1, 
    3606, 
    1, 
    3608, 
    1, 
    3609, 
    1, 
    3610, 
    1, 
    3611, 
    1, 
    3613, 
    1, 
    3614, 
    1, 
    3615, 
    1, 
    3617, 
    1, 
    3617, 
    1, 
    3619, 
    1, 
    3621, 
    1, 
    3622, 
    1, 
    3623, 
    1, 
    3624, 
    1, 
    3626, 
    1, 
    3627, 
    1, 
    3628, 
    1, 
    3630, 
    1, 
    3630, 
    1, 
    3632, 
    1, 
    3634, 
    1, 
    3635, 
    1, 
    3636, 
    1, 
    3637, 
    1, 
    3639, 
    1, 
    3640, 
    1, 
    3641, 
    1, 
    3643, 
    1, 
    3643, 
    1, 
    3645, 
    1, 
    3647, 
    1, 
    3648, 
    1, 
    3649, 
    1, 
    3650, 
    1, 
    3652, 
    1, 
    3653, 
    1, 
    3654, 
    1, 
    3656, 
    1, 
    3656, 
    1, 
    3658, 
    1, 
    3660, 
    1, 
    3661, 
    1, 
    3662, 
    1, 
    3663, 
    1, 
    3665, 
    1, 
    3666, 
    1, 
    3667, 
    1, 
    3669, 
    1, 
    3669, 
    1, 
    3671, 
    1, 
    3673, 
    1, 
    3674, 
    1, 
    3675, 
    1, 
    3676, 
    1, 
    3678, 
    1, 
    3679, 
    1, 
    3680, 
    1, 
    3682, 
    1, 
    3682, 
    1, 
    3684, 
    1, 
    3686, 
    1, 
    3687, 
    1, 
    3688, 
    1, 
    3689, 
    1, 
    3691, 
    1, 
    3692, 
    1, 
    3693, 
    1, 
    3695, 
    1, 
    3695, 
    1, 
    3697, 
    1, 
    3699, 
    1, 
    3699, 
    1, 
    3700, 
    1, 
    3697, 
    1, 
    3694, 
    1, 
    3690, 
    1, 
    3687, 
    1, 
    3684, 
    1, 
    3680, 
    1, 
    3677, 
    1, 
    3674, 
    1, 
    3670, 
    1, 
    3667, 
    1, 
    3664, 
    1, 
    3662, 
    1, 
    3657, 
    1, 
    3655, 
    1, 
    3652, 
    1, 
    3648, 
    1, 
    3645, 
    1, 
    3642, 
    1, 
    3638, 
    1, 
    3635, 
    1, 
    3632, 
    1, 
    3629, 
    1, 
    3625, 
    1, 
    3622, 
    1, 
    3619, 
    1, 
    3615, 
    1, 
    3612, 
    1, 
    3609, 
    1, 
    3605, 
    1, 
    3602, 
    1, 
    3599, 
    1, 
    3596, 
    1, 
    3592, 
    1, 
    3589, 
    1, 
    3586, 
    1, 
    3583, 
    1, 
    3580, 
    1, 
    3577, 
    1, 
    3573, 
    1, 
    3570, 
    1, 
    3567, 
    1, 
    3564, 
    1, 
    3560, 
    1, 
    3557, 
    1, 
    3554, 
    1, 
    3550, 
    1, 
    3547, 
    1, 
    3544, 
    1, 
    3540, 
    1, 
    3537, 
    1, 
    3534, 
    1, 
    3531, 
    1, 
    3527, 
    1, 
    3524, 
    1, 
    3521, 
    1, 
    3517, 
    1, 
    3515, 
    1, 
    3512, 
    1, 
    3508, 
    1, 
    3505, 
    1, 
    3502, 
    1, 
    3499, 
    1, 
    3495, 
    1, 
    3492, 
    1, 
    3489, 
    1, 
    3485, 
    1, 
    3482, 
    1, 
    3479, 
    1, 
    3475, 
    1, 
    3472, 
    1, 
    3469, 
    1, 
    3466, 
    1, 
    3462, 
    1, 
    3461, 
    1, 
    3460, 
    1, 
    3458, 
    1, 
    3457, 
    1, 
    3457, 
    1, 
    3455, 
    1, 
    3454, 
    1, 
    3453, 
    1, 
    3452, 
    1, 
    3450, 
    1, 
    3449, 
    1, 
    3448, 
    1, 
    3447, 
    1, 
    3446, 
    1, 
    3445, 
    1, 
    3443, 
    1, 
    3442, 
    1, 
    3441, 
    1, 
    3440, 
    1, 
    3438, 
    1, 
    3438, 
    1, 
    3437, 
    1, 
    3435, 
    1, 
    3434, 
    1, 
    3433, 
    1, 
    3431, 
    1, 
    3430, 
    1, 
    3429, 
    1, 
    3429, 
    1, 
    3427, 
    1, 
    3426, 
    1, 
    3425, 
    1, 
    3423, 
    1, 
    3422, 
    1, 
    3421, 
    1, 
    3419, 
    1, 
    3419, 
    1, 
    3418, 
    1, 
    3417, 
    1, 
    3415, 
    1, 
    3414, 
    1, 
    3413, 
    1, 
    3411, 
    1, 
    3410, 
    1, 
    3410, 
    1, 
    3408, 
    1, 
    3407, 
    1, 
    3406, 
    1, 
    3405, 
    1, 
    3403, 
    1, 
    3402, 
    1, 
    3401, 
    1, 
    3400, 
    1, 
    3397, 
    1, 
    3393, 
    1, 
    3389, 
    1, 
    3385, 
    1, 
    3381, 
    1, 
    3377, 
    1, 
    3372, 
    1, 
    3369, 
    1, 
    3365, 
    1, 
    3360, 
    1, 
    3356, 
    1, 
    3352, 
    1, 
    3348, 
    1, 
    3344, 
    1, 
    3340, 
    1, 
    3336, 
    1, 
    3331, 
    1, 
    3327, 
    1, 
    3322, 
    1, 
    3317, 
    1, 
    3312, 
    1, 
    3307, 
    1, 
    3302, 
    1, 
    3297, 
    1, 
    3292, 
    1, 
    3288, 
    1, 
    3282, 
    1, 
    3277, 
    1, 
    3273, 
    1, 
    3267, 
    1, 
    3262, 
    1, 
    3258, 
    1, 
    3252, 
    1, 
    3247, 
    1, 
    3243, 
    1, 
    3238, 
    1, 
    3232, 
    1, 
    3229, 
    1, 
    3227, 
    1, 
    3224, 
    1, 
    3221, 
    1, 
    3219, 
    1, 
    3215, 
    1, 
    3213, 
    1, 
    3211, 
    1, 
    3208, 
    1, 
    3205, 
    1, 
    3202, 
    1, 
    3200, 
    1, 
    3197, 
    1, 
    3194, 
    1, 
    3192, 
    1, 
    3188, 
    1, 
    3186, 
    1, 
    3184, 
    1, 
    3181, 
    1, 
    3178, 
    1, 
    3173, 
    1, 
    3169, 
    1, 
    3164, 
    1, 
    3158, 
    1, 
    3154, 
    1, 
    3148, 
    1, 
    3144, 
    1, 
    3139, 
    1, 
    3134, 
    1, 
    3129, 
    1, 
    3125, 
    1, 
    3119, 
    1, 
    3114, 
    1, 
    3109, 
    1, 
    3102, 
    1, 
    3096, 
    1, 
    3089, 
    1, 
    3083, 
    1, 
    3077, 
    1, 
    3071, 
    1, 
    3064, 
    1, 
    3057, 
    1, 
    3052, 
    1, 
    3045, 
    1, 
    3039, 
    1, 
    3032, 
    1, 
    3026, 
    1, 
    3020, 
    1, 
    3014, 
    1, 
    3007, 
    1, 
    3000, 
    1, 
    2995, 
    1, 
    2988, 
    1, 
    2982, 
    1, 
    2975, 
    1, 
    2969, 
    1, 
    2963, 
    1, 
    2957, 
    1, 
    2950, 
    1, 
    2943, 
    1, 
    2938, 
    1, 
    2931, 
    1, 
    2925, 
    1, 
    2917, 
    1, 
    2910, 
    1, 
    2901, 
    1, 
    2894, 
    1, 
    2886, 
    1, 
    2877, 
    1, 
    2870, 
    1, 
    2861, 
    1, 
    2854, 
    1, 
    2845, 
    1, 
    2838, 
    1, 
    2830, 
    1, 
    2822, 
    1, 
    2814, 
    1, 
    2806, 
    1, 
    2798, 
    1, 
    2790, 
    1, 
    2782, 
    1, 
    2774, 
    1, 
    2766, 
    1, 
    2758, 
    1, 
    2750, 
    1, 
    2742, 
    1, 
    2735, 
    1, 
    2726, 
    1, 
    2718, 
    1, 
    2710, 
    1, 
    2702, 
    1, 
    2694, 
    1, 
    2686, 
    1, 
    2679, 
    1, 
    2670, 
    1, 
    2663, 
    1, 
    2654, 
    1, 
    2646, 
    1, 
    2639, 
    1, 
    2630, 
    1, 
    2623, 
    1, 
    2614, 
    1, 
    2607, 
    1, 
    2598, 
    1, 
    2591, 
    1, 
    2582, 
    1, 
    2574, 
    1, 
    2567, 
    1, 
    2558, 
    1, 
    2551, 
    1, 
    2542, 
    1, 
    2535, 
    1, 
    2527, 
    1, 
    2519, 
    1, 
    2511, 
    1, 
    2502, 
    1, 
    2495, 
    1, 
    2486, 
    1, 
    2479, 
    1, 
    2471, 
    1, 
    2463, 
    1, 
    2455, 
    1, 
    2447, 
    1, 
    2439, 
    1, 
    2430, 
    1, 
    2423, 
    1, 
    2415, 
    1, 
    2407, 
    1, 
    2399, 
    1, 
    2391, 
    1, 
    2383, 
    1, 
    2375, 
    1, 
    2367, 
    1, 
    2359, 
    1, 
    2351, 
    1, 
    2343, 
    1, 
    2335, 
    1, 
    2327, 
    1, 
    2320, 
    1, 
    2311, 
    1, 
    2304, 
    1, 
    2295, 
    1, 
    2287, 
    1, 
    2279, 
    1, 
    2271, 
    1, 
    2263, 
    1, 
    2255, 
    1, 
    2248, 
    1, 
    2239, 
    1, 
    2232, 
    1, 
    2223, 
    1, 
    2215, 
    1, 
    2208, 
    1, 
    2199, 
    1, 
    2192, 
    1, 
    2183, 
    1, 
    2176, 
    1, 
    2167, 
    1, 
    2160, 
    1, 
    2152, 
    1, 
    2143, 
    1, 
    2136, 
    1, 
    2127, 
    1, 
    2120, 
    1, 
    2111, 
    1, 
    2104, 
    1, 
    2096, 
    1, 
    2088, 
    1, 
    2080, 
    1, 
    2072, 
    1, 
    2064, 
    1, 
    2055, 
    1, 
    2048, 
    1, 
    2040, 
    1, 
    2032, 
    1, 
    2024, 
    1, 
    2016, 
    1, 
    2008, 
    1, 
    2001, 
    1, 
    1992, 
    1, 
    1984, 
    1, 
    1976, 
    1, 
    1968, 
    1, 
    1960, 
    1, 
    1952, 
    1, 
    1945, 
    1, 
    1936, 
    1, 
    1929, 
    1, 
    1920, 
    1, 
    1912, 
    1, 
    1904, 
    1, 
    1896, 
    1, 
    1889, 
    1, 
    1880, 
    1, 
    1873, 
    1, 
    1864, 
    1, 
    1857, 
    1, 
    1848, 
    1, 
    1840, 
    1, 
    1833, 
    1, 
    1824, 
    1, 
    1817, 
    1, 
    1808, 
    1, 
    1801, 
    1, 
    1792, 
    1, 
    1785, 
    1, 
    1777, 
    1, 
    1768, 
    1, 
    1761, 
    1, 
    1752, 
    1, 
    1745, 
    1, 
    1736, 
    1, 
    1729, 
    1, 
    1721, 
    1, 
    1713, 
    1, 
    1705, 
    1, 
    1696, 
    1, 
    1689, 
    1, 
    1681, 
    1, 
    1673, 
    1, 
    1665, 
    1, 
    1657, 
    1, 
    1649, 
    1, 
    1641, 
    1, 
    1633, 
    1, 
    1625, 
    1, 
    1617, 
    1, 
    1609, 
    1, 
    1601, 
    1, 
    1593, 
    1, 
    1585, 
    1, 
    1577, 
    1, 
    1570, 
    1, 
    1561, 
    1, 
    1553, 
    1, 
    1545, 
    1, 
    1537, 
    1, 
    1529, 
    1, 
    1521, 
    1, 
    1514, 
    1, 
    1505, 
    1, 
    1498, 
    1, 
    1489, 
    1, 
    1481, 
    1, 
    1473, 
    1, 
    1465, 
    1, 
    1458, 
    1, 
    1449, 
    1, 
    1442, 
    1, 
    1433, 
    1, 
    1426, 
    1, 
    1417, 
    1, 
    1409, 
    1, 
    1402, 
    1, 
    1393, 
    1, 
    1386, 
    1, 
    1377, 
    1, 
    1370, 
    1, 
    1362, 
    1, 
    1354, 
    1, 
    1346, 
    1, 
    1338, 
    1, 
    1330, 
    1, 
    1321, 
    1, 
    1314, 
    1, 
    1306, 
    1, 
    1298, 
    1, 
    1290, 
    1, 
    1282, 
    1, 
    1274, 
    1, 
    1266, 
    1, 
    1258, 
    1, 
    1250, 
    1, 
    1242, 
    1, 
    1234, 
    1, 
    1226, 
    1, 
    1218, 
    1, 
    1210, 
    1, 
    1202, 
    1, 
    1195, 
    1, 
    1186, 
    1, 
    1178, 
    1, 
    1170, 
    1, 
    1162, 
    1, 
    1154, 
    1, 
    1146, 
    1, 
    1139, 
    1, 
    1130, 
    1, 
    1123, 
    1, 
    1114, 
    1, 
    1106, 
    1, 
    1098, 
    1, 
    1090, 
    1, 
    1083, 
    1, 
    1074, 
    1, 
    1067, 
    1, 
    1058, 
    1, 
    1051, 
    1, 
    1043, 
    1, 
    1034, 
    1, 
    1027, 
    1, 
    1018, 
    1, 
    1011, 
    1, 
    1002, 
    1, 
    995, 
    1, 
    987, 
    1, 
    971, 
    1, 
    923, 
    1, 
    872, 
    1, 
    825, 
    1, 
    775, 
    1, 
    727, 
    1, 
    676, 
    1, 
    629, 
    1, 
    579, 
    1, 
    530, 
    1, 
    480, 
    1, 
    432, 
    1, 
    383, 
    1, 
    333, 
    1, 
    285, 
    1, 
    236, 
    1, 
    187, 
    1, 
    137, 
    1, 
    89, 
    1, 40 ;

 runvals = 
    188381733, 
    21599, 
    1, 
    21597, 
    1, 
    21594, 
    1, 
    21592, 
    1, 
    21590, 
    1, 
    21588, 
    1, 
    21585, 
    1, 
    21583, 
    1, 
    21581, 
    1, 
    21579, 
    1, 
    21575, 
    1, 
    21573, 
    1, 
    21571, 
    1, 
    21569, 
    1, 
    21566, 
    1, 
    21564, 
    1, 
    21562, 
    1, 
    21560, 
    1, 
    21557, 
    1, 
    21555, 
    1, 
    21553, 
    1, 
    21551, 
    1, 
    21548, 
    1, 
    21546, 
    1, 
    21544, 
    1, 
    21541, 
    1, 
    21539, 
    1, 
    21537, 
    1, 
    21535, 
    1, 
    21532, 
    1, 
    21530, 
    1, 
    21528, 
    1, 
    21526, 
    1, 
    21523, 
    1, 
    21521, 
    1, 
    21519, 
    1, 
    21517, 
    1, 
    21514, 
    1, 
    21512, 
    1, 
    21510, 
    1, 
    21507, 
    1, 
    21504, 
    1, 
    21502, 
    1, 
    21500, 
    1, 
    21498, 
    1, 
    21495, 
    1, 
    21493, 
    1, 
    21491, 
    1, 
    21489, 
    1, 
    21486, 
    1, 
    21484, 
    1, 
    21482, 
    1, 
    21479, 
    1, 
    21477, 
    1, 
    21475, 
    1, 
    21473, 
    1, 
    21470, 
    1, 
    21468, 
    1, 
    21466, 
    1, 
    21464, 
    1, 
    21461, 
    1, 
    21459, 
    1, 
    21457, 
    1, 
    21455, 
    1, 
    21452, 
    1, 
    21450, 
    1, 
    21448, 
    1, 
    21446, 
    1, 
    21443, 
    1, 
    21441, 
    1, 
    21438, 
    1, 
    21436, 
    1, 
    21433, 
    1, 
    21431, 
    1, 
    21429, 
    1, 
    21426, 
    1, 
    21424, 
    1, 
    21422, 
    1, 
    21420, 
    1, 
    21417, 
    1, 
    21415, 
    1, 
    21413, 
    1, 
    21411, 
    1, 
    21408, 
    1, 
    21406, 
    1, 
    21404, 
    1, 
    21402, 
    1, 
    21399, 
    1, 
    21397, 
    1, 
    21395, 
    1, 
    21393, 
    1, 
    21390, 
    1, 
    21388, 
    1, 
    21386, 
    1, 
    21384, 
    1, 
    21381, 
    1, 
    21379, 
    1, 
    21377, 
    1, 
    21375, 
    1, 
    21372, 
    1, 
    21370, 
    1, 
    21367, 
    1, 
    21364, 
    1, 
    21362, 
    1, 
    21360, 
    1, 
    21358, 
    1, 
    21355, 
    1, 
    21353, 
    1, 
    21351, 
    1, 
    21349, 
    1, 
    21346, 
    1, 
    21344, 
    1, 
    21342, 
    1, 
    21340, 
    1, 
    21337, 
    1, 
    21335, 
    1, 
    21333, 
    1, 
    21331, 
    1, 
    21328, 
    1, 
    21326, 
    1, 
    21324, 
    1, 
    21322, 
    1, 
    21319, 
    1, 
    21317, 
    1, 
    21315, 
    1, 
    21312, 
    1, 
    21310, 
    1, 
    21308, 
    1, 
    21306, 
    1, 
    21303, 
    1, 
    21301, 
    1, 
    21298, 
    1, 
    21296, 
    1, 
    21293, 
    1, 
    21291, 
    1, 
    21289, 
    1, 
    21287, 
    1, 
    21284, 
    1, 
    21282, 
    1, 
    21280, 
    1, 
    21278, 
    1, 
    21275, 
    1, 
    21273, 
    1, 
    21271, 
    1, 
    21269, 
    1, 
    21266, 
    1, 
    21264, 
    1, 
    21262, 
    1, 
    21260, 
    1, 
    21257, 
    1, 
    21255, 
    1, 
    21253, 
    1, 
    21250, 
    1, 
    21248, 
    1, 
    21246, 
    1, 
    21244, 
    1, 
    21241, 
    1, 
    21239, 
    1, 
    21237, 
    1, 
    21235, 
    1, 
    21232, 
    1, 
    21230, 
    1, 
    21227, 
    1, 
    21225, 
    1, 
    21222, 
    1, 
    21220, 
    1, 
    21218, 
    1, 
    21216, 
    1, 
    21213, 
    1, 
    21211, 
    1, 
    21209, 
    1, 
    21207, 
    1, 
    21204, 
    1, 
    21202, 
    1, 
    21200, 
    1, 
    21197, 
    1, 
    21195, 
    1, 
    21193, 
    1, 
    21191, 
    1, 
    21188, 
    1, 
    21186, 
    1, 
    21184, 
    1, 
    21182, 
    1, 
    21179, 
    1, 
    21177, 
    1, 
    21175, 
    1, 
    21173, 
    1, 
    21170, 
    1, 
    21168, 
    1, 
    21166, 
    1, 
    21164, 
    1, 
    21161, 
    1, 
    21158, 
    1, 
    21156, 
    1, 
    21154, 
    1, 
    21151, 
    1, 
    21149, 
    1, 
    21147, 
    1, 
    21145, 
    1, 
    21142, 
    1, 
    21140, 
    1, 
    21138, 
    1, 
    21135, 
    1, 
    21133, 
    1, 
    21131, 
    1, 
    21129, 
    1, 
    21126, 
    1, 
    21124, 
    1, 
    21122, 
    1, 
    21120, 
    1, 
    21117, 
    1, 
    21115, 
    1, 
    21113, 
    1, 
    21111, 
    1, 
    21108, 
    1, 
    21106, 
    1, 
    21104, 
    1, 
    21102, 
    1, 
    21099, 
    1, 
    21097, 
    1, 
    21095, 
    1, 
    21093, 
    1, 
    21089, 
    1, 
    21087, 
    1, 
    21085, 
    1, 
    21082, 
    1, 
    21080, 
    1, 
    21078, 
    1, 
    21076, 
    1, 
    21073, 
    1, 
    21071, 
    1, 
    21069, 
    1, 
    21067, 
    1, 
    21064, 
    1, 
    21062, 
    1, 
    21060, 
    1, 
    21058, 
    1, 
    21055, 
    1, 
    21053, 
    1, 
    21051, 
    1, 
    21049, 
    1, 
    21046, 
    1, 
    21044, 
    1, 
    21042, 
    1, 
    21040, 
    1, 
    21037, 
    1, 
    21035, 
    1, 
    21033, 
    1, 
    21031, 
    1, 
    21028, 
    1, 
    21026, 
    1, 
    21024, 
    1, 
    21020, 
    1, 
    21018, 
    1, 
    21016, 
    1, 
    21014, 
    1, 
    21011, 
    1, 
    21009, 
    1, 
    21007, 
    1, 
    21005, 
    1, 
    21002, 
    1, 
    21000, 
    1, 
    20998, 
    1, 
    20996, 
    1, 
    20993, 
    1, 
    20991, 
    1, 
    20989, 
    1, 
    20987, 
    1, 
    20984, 
    1, 
    20982, 
    1, 
    20980, 
    1, 
    20978, 
    1, 
    20975, 
    1, 
    20973, 
    1, 
    20971, 
    1, 
    20968, 
    1, 
    20966, 
    1, 
    20964, 
    1, 
    20962, 
    1, 
    20959, 
    1, 
    20957, 
    1, 
    20955, 
    1, 
    20953, 
    1, 
    20949, 
    1, 
    20947, 
    1, 
    20945, 
    1, 
    20943, 
    1, 
    20940, 
    1, 
    20938, 
    1, 
    20936, 
    1, 
    20934, 
    1, 
    20931, 
    1, 
    20929, 
    1, 
    20927, 
    1, 
    20925, 
    1, 
    20922, 
    1, 
    20920, 
    1, 
    20918, 
    1, 
    20916, 
    1, 
    20913, 
    1, 
    20911, 
    1, 
    20909, 
    1, 
    20906, 
    1, 
    20904, 
    1, 
    20902, 
    1, 
    20900, 
    1, 
    20897, 
    1, 
    20895, 
    1, 
    20893, 
    1, 
    20891, 
    1, 
    20888, 
    1, 
    20886, 
    1, 
    20884, 
    1, 
    20882, 
    1, 
    20878, 
    1, 
    20876, 
    1, 
    20874, 
    1, 
    20872, 
    1, 
    20869, 
    1, 
    20867, 
    1, 
    20865, 
    1, 
    20863, 
    1, 
    20860, 
    1, 
    20858, 
    1, 
    20856, 
    1, 
    20853, 
    1, 
    20851, 
    1, 
    20849, 
    1, 
    20847, 
    1, 
    20844, 
    1, 
    20842, 
    1, 
    20840, 
    1, 
    20838, 
    1, 
    20835, 
    1, 
    20833, 
    1, 
    20831, 
    1, 
    20829, 
    1, 
    20826, 
    1, 
    20824, 
    1, 
    20822, 
    1, 
    20820, 
    1, 
    20817, 
    1, 
    20815, 
    1, 
    20813, 
    1, 
    20810, 
    1, 
    20807, 
    1, 
    20805, 
    1, 
    20803, 
    1, 
    20801, 
    1, 
    20798, 
    1, 
    20796, 
    1, 
    20794, 
    1, 
    20791, 
    1, 
    20789, 
    1, 
    20787, 
    1, 
    20785, 
    1, 
    20782, 
    1, 
    20780, 
    1, 
    20778, 
    1, 
    20776, 
    1, 
    20773, 
    1, 
    20771, 
    1, 
    20769, 
    1, 
    20767, 
    1, 
    20764, 
    1, 
    20762, 
    1, 
    20760, 
    1, 
    20758, 
    1, 
    20755, 
    1, 
    20753, 
    1, 
    20751, 
    1, 
    20749, 
    1, 
    20746, 
    1, 
    20744, 
    1, 
    20741, 
    1, 
    20738, 
    1, 
    20736, 
    1, 
    20734, 
    1, 
    20732, 
    1, 
    20729, 
    1, 
    20727, 
    1, 
    20725, 
    1, 
    20723, 
    1, 
    20720, 
    1, 
    20718, 
    1, 
    20716, 
    1, 
    20714, 
    1, 
    20711, 
    1, 
    20709, 
    1, 
    20707, 
    1, 
    20705, 
    1, 
    20702, 
    1, 
    20700, 
    1, 
    20698, 
    1, 
    20696, 
    1, 
    20693, 
    1, 
    20691, 
    1, 
    20689, 
    1, 
    20687, 
    1, 
    20684, 
    1, 
    20682, 
    1, 
    20680, 
    1, 
    20678, 
    1, 
    20675, 
    1, 
    20673, 
    1, 
    20670, 
    1, 
    20667, 
    1, 
    20665, 
    1, 
    20663, 
    1, 
    20661, 
    1, 
    20658, 
    1, 
    20656, 
    1, 
    20654, 
    1, 
    20652, 
    1, 
    20649, 
    1, 
    20647, 
    1, 
    20645, 
    1, 
    20643, 
    1, 
    20640, 
    1, 
    20638, 
    1, 
    20636, 
    1, 
    20634, 
    1, 
    20631, 
    1, 
    20629, 
    1, 
    20627, 
    1, 
    20624, 
    1, 
    20622, 
    1, 
    20620, 
    1, 
    20618, 
    1, 
    20615, 
    1, 
    20613, 
    1, 
    20611, 
    1, 
    20609, 
    1, 
    20606, 
    1, 
    20604, 
    1, 
    20601, 
    1, 
    20599, 
    1, 
    20596, 
    1, 
    20594, 
    1, 
    20592, 
    1, 
    20590, 
    1, 
    20587, 
    1, 
    20585, 
    1, 
    20583, 
    1, 
    20581, 
    1, 
    20578, 
    1, 
    20576, 
    1, 
    20574, 
    1, 
    20572, 
    1, 
    20569, 
    1, 
    20567, 
    1, 
    20565, 
    1, 
    20563, 
    1, 
    20560, 
    1, 
    20558, 
    1, 
    20556, 
    1, 
    20553, 
    1, 
    20551, 
    1, 
    20549, 
    1, 
    20547, 
    1, 
    20544, 
    1, 
    20542, 
    1, 
    20540, 
    1, 
    20538, 
    1, 
    20535, 
    1, 
    20533, 
    1, 
    20530, 
    1, 
    20528, 
    1, 
    20525, 
    1, 
    20523, 
    1, 
    20521, 
    1, 
    20519, 
    1, 
    20516, 
    1, 
    20514, 
    1, 
    20512, 
    1, 
    20509, 
    1, 
    20507, 
    1, 
    20505, 
    1, 
    20503, 
    1, 
    20500, 
    1, 
    20498, 
    1, 
    20496, 
    1, 
    20494, 
    1, 
    20491, 
    1, 
    20489, 
    1, 
    20487, 
    1, 
    20485, 
    1, 
    20482, 
    1, 
    20480, 
    1, 
    20478, 
    1, 
    20476, 
    1, 
    20473, 
    1, 
    20471, 
    1, 
    20469, 
    1, 
    20467, 
    1, 
    20464, 
    1, 
    20461, 
    1, 
    20459, 
    1, 
    20457, 
    1, 
    20454, 
    1, 
    20452, 
    1, 
    20450, 
    1, 
    20447, 
    1, 
    20445, 
    1, 
    20443, 
    1, 
    20441, 
    1, 
    20438, 
    1, 
    20436, 
    1, 
    20434, 
    1, 
    20432, 
    1, 
    20429, 
    1, 
    20427, 
    1, 
    20425, 
    1, 
    20423, 
    1, 
    20420, 
    1, 
    20418, 
    1, 
    20416, 
    1, 
    20414, 
    1, 
    20411, 
    1, 
    20409, 
    1, 
    20407, 
    1, 
    20405, 
    1, 
    20402, 
    1, 
    20400, 
    1, 
    20398, 
    1, 
    20395, 
    1, 
    20392, 
    1, 
    20390, 
    1, 
    20388, 
    1, 
    20385, 
    1, 
    20383, 
    1, 
    20381, 
    1, 
    20379, 
    1, 
    20376, 
    1, 
    20374, 
    1, 
    20372, 
    1, 
    20370, 
    1, 
    20367, 
    1, 
    20365, 
    1, 
    20363, 
    1, 
    20361, 
    1, 
    20358, 
    1, 
    20356, 
    1, 
    20354, 
    1, 
    20352, 
    1, 
    20349, 
    1, 
    20347, 
    1, 
    20345, 
    1, 
    20343, 
    1, 
    20340, 
    1, 
    20338, 
    1, 
    20336, 
    1, 
    20333, 
    1, 
    20331, 
    1, 
    20329, 
    1, 
    20327, 
    1, 
    20324, 
    1, 
    20321, 
    1, 
    20319, 
    1, 
    20317, 
    1, 
    20314, 
    1, 
    20312, 
    1, 
    20310, 
    1, 
    20308, 
    1, 
    20305, 
    1, 
    20303, 
    1, 
    20301, 
    1, 
    20299, 
    1, 
    20296, 
    1, 
    20294, 
    1, 
    20292, 
    1, 
    20290, 
    1, 
    20287, 
    1, 
    20285, 
    1, 
    20283, 
    1, 
    20280, 
    1, 
    20278, 
    1, 
    20276, 
    1, 
    20274, 
    1, 
    20271, 
    1, 
    20269, 
    1, 
    20267, 
    1, 
    20265, 
    1, 
    20262, 
    1, 
    20260, 
    1, 
    20258, 
    1, 
    20256, 
    1, 
    20252, 
    1, 
    20250, 
    1, 
    20248, 
    1, 
    20246, 
    1, 
    20243, 
    1, 
    20241, 
    1, 
    20239, 
    1, 
    20237, 
    1, 
    20234, 
    1, 
    20232, 
    1, 
    20230, 
    1, 
    20228, 
    1, 
    20225, 
    1, 
    20223, 
    1, 
    20221, 
    1, 
    20218, 
    1, 
    20216, 
    1, 
    20214, 
    1, 
    20212, 
    1, 
    20209, 
    1, 
    20207, 
    1, 
    20205, 
    1, 
    20203, 
    1, 
    20200, 
    1, 
    20198, 
    1, 
    20196, 
    1, 
    20194, 
    1, 
    20191, 
    1, 
    20189, 
    1, 
    20187, 
    1, 
    20185, 
    1, 
    20181, 
    1, 
    20179, 
    1, 
    20177, 
    1, 
    20175, 
    1, 
    20172, 
    1, 
    20170, 
    1, 
    20168, 
    1, 
    20165, 
    1, 
    20163, 
    1, 
    20161, 
    1, 
    20159, 
    1, 
    20156, 
    1, 
    20154, 
    1, 
    20152, 
    1, 
    20150, 
    1, 
    20147, 
    1, 
    20145, 
    1, 
    20143, 
    1, 
    20141, 
    1, 
    20138, 
    1, 
    20136, 
    1, 
    20134, 
    1, 
    20132, 
    1, 
    20129, 
    1, 
    20127, 
    1, 
    20125, 
    1, 
    20123, 
    1, 
    20120, 
    1, 
    20118, 
    1, 
    20116, 
    1, 
    20113, 
    1, 
    20110, 
    1, 
    20108, 
    1, 
    20106, 
    1, 
    20103, 
    1, 
    20101, 
    1, 
    20099, 
    1, 
    20097, 
    1, 
    20094, 
    1, 
    20092, 
    1, 
    20090, 
    1, 
    20088, 
    1, 
    20085, 
    1, 
    20083, 
    1, 
    20081, 
    1, 
    20079, 
    1, 
    20076, 
    1, 
    20074, 
    1, 
    20072, 
    1, 
    20068, 
    1, 
    20063, 
    1, 
    20058, 
    1, 
    20054, 
    1, 
    20049, 
    1, 
    20045, 
    1, 
    20040, 
    1, 
    20036, 
    1, 
    20031, 
    1, 
    20026, 
    1, 
    20022, 
    1, 
    20016, 
    1, 
    20012, 
    1, 
    20007, 
    1, 
    20003, 
    1, 
    19998, 
    1, 
    19993, 
    1, 
    19989, 
    1, 
    19984, 
    1, 
    19980, 
    1, 
    19975, 
    1, 
    19971, 
    1, 
    19966, 
    1, 
    19962, 
    1, 
    19957, 
    1, 
    19952, 
    1, 
    19948, 
    1, 
    19943, 
    1, 
    19939, 
    1, 
    19934, 
    1, 
    19930, 
    1, 
    19925, 
    1, 
    19920, 
    1, 
    19916, 
    1, 
    19911, 
    1, 
    19907, 
    1, 
    19902, 
    1, 
    19898, 
    1, 
    19893, 
    1, 
    19888, 
    1, 
    19884, 
    1, 
    19879, 
    1, 
    19874, 
    1, 
    19869, 
    1, 
    19865, 
    1, 
    19860, 
    1, 
    19855, 
    1, 
    19851, 
    1, 
    19846, 
    1, 
    19842, 
    1, 
    19837, 
    1, 
    19833, 
    1, 
    19828, 
    1, 
    19824, 
    1, 
    19819, 
    1, 
    19814, 
    1, 
    19810, 
    1, 
    19805, 
    1, 
    19801, 
    1, 
    19796, 
    1, 
    19792, 
    1, 
    19787, 
    1, 
    19782, 
    1, 
    19778, 
    1, 
    19773, 
    1, 
    19769, 
    1, 
    19764, 
    1, 
    19760, 
    1, 
    19755, 
    1, 
    19750, 
    1, 
    19746, 
    1, 
    19741, 
    1, 
    19736, 
    1, 
    19731, 
    1, 
    19727, 
    1, 
    19722, 
    1, 
    19717, 
    1, 
    19713, 
    1, 
    19708, 
    1, 
    19704, 
    1, 
    19699, 
    1, 
    19695, 
    1, 
    19690, 
    1, 
    19686, 
    1, 
    19681, 
    1, 
    19677, 
    1, 
    19672, 
    1, 
    19667, 
    1, 
    19663, 
    1, 
    19658, 
    1, 
    19654, 
    1, 
    19649, 
    1, 
    19644, 
    1, 
    19640, 
    1, 
    19635, 
    1, 
    19631, 
    1, 
    19626, 
    1, 
    19622, 
    1, 
    19617, 
    1, 
    19612, 
    1, 
    19608, 
    1, 
    19603, 
    1, 
    19599, 
    1, 
    19593, 
    1, 
    19589, 
    1, 
    19584, 
    1, 
    19579, 
    1, 
    19575, 
    1, 
    19570, 
    1, 
    19566, 
    1, 
    19561, 
    1, 
    19557, 
    1, 
    19552, 
    1, 
    19548, 
    1, 
    19543, 
    1, 
    19538, 
    1, 
    19534, 
    1, 
    19529, 
    1, 
    19525, 
    1, 
    19520, 
    1, 
    19516, 
    1, 
    19511, 
    1, 
    19506, 
    1, 
    19502, 
    1, 
    19497, 
    1, 
    19493, 
    1, 
    19488, 
    1, 
    19484, 
    1, 
    19479, 
    1, 
    19474, 
    1, 
    19470, 
    1, 
    19465, 
    1, 
    19461, 
    1, 
    19455, 
    1, 
    19451, 
    1, 
    19446, 
    1, 
    19441, 
    1, 
    19437, 
    1, 
    19432, 
    1, 
    19428, 
    1, 
    19423, 
    1, 
    19419, 
    1, 
    19414, 
    1, 
    19410, 
    1, 
    19405, 
    1, 
    19400, 
    1, 
    19396, 
    1, 
    19391, 
    1, 
    19387, 
    1, 
    19382, 
    1, 
    19378, 
    1, 
    19373, 
    1, 
    19368, 
    1, 
    19364, 
    1, 
    19359, 
    1, 
    19355, 
    1, 
    19350, 
    1, 
    19346, 
    1, 
    19341, 
    1, 
    19336, 
    1, 
    19332, 
    1, 
    19327, 
    1, 
    19323, 
    1, 
    19317, 
    1, 
    19313, 
    1, 
    19308, 
    1, 
    19303, 
    1, 
    19299, 
    1, 
    19294, 
    1, 
    19290, 
    1, 
    19285, 
    1, 
    19281, 
    1, 
    19276, 
    1, 
    19272, 
    1, 
    19267, 
    1, 
    19263, 
    1, 
    19258, 
    1, 
    19253, 
    1, 
    19249, 
    1, 
    19244, 
    1, 
    19240, 
    1, 
    19235, 
    1, 
    19230, 
    1, 
    19226, 
    1, 
    19221, 
    1, 
    19217, 
    1, 
    19212, 
    1, 
    19208, 
    1, 
    19203, 
    1, 
    19198, 
    1, 
    19194, 
    1, 
    19189, 
    1, 
    19185, 
    1, 
    19180, 
    1, 
    19175, 
    1, 
    19170, 
    1, 
    19165, 
    1, 
    19161, 
    1, 
    19156, 
    1, 
    19152, 
    1, 
    19150, 
    1, 
    19148, 
    1, 
    19146, 
    1, 
    19145, 
    1, 
    19143, 
    1, 
    19141, 
    1, 
    19140, 
    1, 
    19138, 
    1, 
    19136, 
    1, 
    19134, 
    1, 
    19133, 
    1, 
    19131, 
    1, 
    19129, 
    1, 
    19128, 
    1, 
    19126, 
    1, 
    19124, 
    1, 
    19123, 
    1, 
    19121, 
    1, 
    19119, 
    1, 
    19117, 
    1, 
    19116, 
    1, 
    19114, 
    1, 
    19112, 
    1, 
    19111, 
    1, 
    19108, 
    1, 
    19106, 
    1, 
    19105, 
    1, 
    19103, 
    1, 
    19101, 
    1, 
    19099, 
    1, 
    19098, 
    1, 
    19096, 
    1, 
    19094, 
    1, 
    19093, 
    1, 
    19091, 
    1, 
    19089, 
    1, 
    19088, 
    1, 
    19086, 
    1, 
    19084, 
    1, 
    19082, 
    1, 
    19081, 
    1, 
    19079, 
    1, 
    19077, 
    1, 
    19076, 
    1, 
    19074, 
    1, 
    19072, 
    1, 
    19071, 
    1, 
    19069, 
    1, 
    19067, 
    1, 
    19065, 
    1, 
    19064, 
    1, 
    19062, 
    1, 
    19060, 
    1, 
    19059, 
    1, 
    19057, 
    1, 
    19054, 
    1, 
    19053, 
    1, 
    19051, 
    1, 
    19049, 
    1, 
    19047, 
    1, 
    19046, 
    1, 
    19044, 
    1, 
    19042, 
    1, 
    19041, 
    1, 
    19039, 
    1, 
    19037, 
    1, 
    19036, 
    1, 
    19034, 
    1, 
    19032, 
    1, 
    19030, 
    1, 
    19029, 
    1, 
    19027, 
    1, 
    19025, 
    1, 
    19024, 
    1, 
    19022, 
    1, 
    19020, 
    1, 
    19019, 
    1, 
    19017, 
    1, 
    19015, 
    1, 
    19013, 
    1, 
    19012, 
    1, 
    19010, 
    1, 
    19008, 
    1, 
    19007, 
    1, 
    19005, 
    1, 
    19002, 
    1, 
    19001, 
    1, 
    18999, 
    1, 
    18997, 
    1, 
    18995, 
    1, 
    18994, 
    1, 
    18992, 
    1, 
    18990, 
    1, 
    18989, 
    1, 
    18987, 
    1, 
    18985, 
    1, 
    18984, 
    1, 
    18982, 
    1, 
    18980, 
    1, 
    18979, 
    1, 
    18977, 
    1, 
    18975, 
    1, 
    18973, 
    1, 
    18972, 
    1, 
    18970, 
    1, 
    18968, 
    1, 
    18967, 
    1, 
    18965, 
    1, 
    18963, 
    1, 
    18962, 
    1, 
    18960, 
    1, 
    18958, 
    1, 
    18956, 
    1, 
    18955, 
    1, 
    18953, 
    1, 
    18950, 
    1, 
    18949, 
    1, 
    18947, 
    1, 
    18945, 
    1, 
    18944, 
    1, 
    18942, 
    1, 
    18940, 
    1, 
    18938, 
    1, 
    18937, 
    1, 
    18935, 
    1, 
    18933, 
    1, 
    18932, 
    1, 
    18930, 
    1, 
    18928, 
    1, 
    18927, 
    1, 
    18925, 
    1, 
    18923, 
    1, 
    18921, 
    1, 
    18920, 
    1, 
    18918, 
    1, 
    18916, 
    1, 
    18915, 
    1, 
    18913, 
    1, 
    18911, 
    1, 
    18910, 
    1, 
    18908, 
    1, 
    18906, 
    1, 
    18904, 
    1, 
    18903, 
    1, 
    18901, 
    1, 
    18898, 
    1, 
    18895, 
    1, 
    18892, 
    1, 
    18888, 
    1, 
    18885, 
    1, 
    18881, 
    1, 
    18877, 
    1, 
    18874, 
    1, 
    18871, 
    1, 
    18867, 
    1, 
    18863, 
    1, 
    18860, 
    1, 
    18857, 
    1, 
    18853, 
    1, 
    18850, 
    1, 
    18846, 
    1, 
    18842, 
    1, 
    18839, 
    1, 
    18836, 
    1, 
    18832, 
    1, 
    18828, 
    1, 
    18825, 
    1, 
    18822, 
    1, 
    18818, 
    1, 
    18815, 
    1, 
    18811, 
    1, 
    18808, 
    1, 
    18804, 
    1, 
    18801, 
    1, 
    18797, 
    1, 
    18793, 
    1, 
    18791, 
    1, 
    18787, 
    1, 
    18783, 
    1, 
    18780, 
    1, 
    18776, 
    1, 
    18773, 
    1, 
    18769, 
    1, 
    18766, 
    1, 
    18762, 
    1, 
    18758, 
    1, 
    18756, 
    1, 
    18752, 
    1, 
    18748, 
    1, 
    18745, 
    1, 
    18741, 
    1, 
    18738, 
    1, 
    18734, 
    1, 
    18731, 
    1, 
    18727, 
    1, 
    18723, 
    1, 
    18721, 
    1, 
    18717, 
    1, 
    18713, 
    1, 
    18710, 
    1, 
    18706, 
    1, 
    18703, 
    1, 
    18699, 
    1, 
    18696, 
    1, 
    18692, 
    1, 
    18688, 
    1, 
    18686, 
    1, 
    18682, 
    1, 
    18678, 
    1, 
    18675, 
    1, 
    18671, 
    1, 
    18668, 
    1, 
    18664, 
    1, 
    18661, 
    1, 
    18657, 
    1, 
    18653, 
    1, 
    18651, 
    1, 
    18647, 
    1, 
    18643, 
    1, 
    18640, 
    1, 
    18636, 
    1, 
    18633, 
    1, 
    18629, 
    1, 
    18626, 
    1, 
    18622, 
    1, 
    18618, 
    1, 
    18616, 
    1, 
    18612, 
    1, 
    18608, 
    1, 
    18605, 
    1, 
    18601, 
    1, 
    18598, 
    1, 
    18594, 
    1, 
    18591, 
    1, 
    18587, 
    1, 
    18583, 
    1, 
    18581, 
    1, 
    18577, 
    1, 
    18573, 
    1, 
    18570, 
    1, 
    18567, 
    1, 
    18563, 
    1, 
    18559, 
    1, 
    18556, 
    1, 
    18552, 
    1, 
    18549, 
    1, 
    18546, 
    1, 
    18542, 
    1, 
    18538, 
    1, 
    18535, 
    1, 
    18532, 
    1, 
    18528, 
    1, 
    18524, 
    1, 
    18521, 
    1, 
    18517, 
    1, 
    18514, 
    1, 
    18511, 
    1, 
    18507, 
    1, 
    18503, 
    1, 
    18500, 
    1, 
    18497, 
    1, 
    18493, 
    1, 
    18489, 
    1, 
    18486, 
    1, 
    18482, 
    1, 
    18479, 
    1, 
    18476, 
    1, 
    18472, 
    1, 
    18468, 
    1, 
    18465, 
    1, 
    18462, 
    1, 
    18458, 
    1, 
    18454, 
    1, 
    18451, 
    1, 
    18447, 
    1, 
    18444, 
    1, 
    18441, 
    1, 
    18437, 
    1, 
    18433, 
    1, 
    18430, 
    1, 
    18427, 
    1, 
    18423, 
    1, 
    18419, 
    1, 
    18416, 
    1, 
    18412, 
    1, 
    18409, 
    1, 
    18406, 
    1, 
    18402, 
    1, 
    18398, 
    1, 
    18395, 
    1, 
    18392, 
    1, 
    18388, 
    1, 
    18384, 
    1, 
    18381, 
    1, 
    18377, 
    1, 
    18374, 
    1, 
    18371, 
    1, 
    18367, 
    1, 
    18363, 
    1, 
    18360, 
    1, 
    18357, 
    1, 
    18353, 
    1, 
    18349, 
    1, 
    18346, 
    1, 
    18342, 
    1, 
    18339, 
    1, 
    18336, 
    1, 
    18332, 
    1, 
    18328, 
    1, 
    18326, 
    1, 
    18322, 
    1, 
    18318, 
    1, 
    18315, 
    1, 
    18311, 
    1, 
    18308, 
    1, 
    18304, 
    1, 
    18301, 
    1, 
    18297, 
    1, 
    18293, 
    1, 
    18291, 
    1, 
    18287, 
    1, 
    18283, 
    1, 
    18280, 
    1, 
    18276, 
    1, 
    18273, 
    1, 
    18269, 
    1, 
    18266, 
    1, 
    18262, 
    1, 
    18258, 
    1, 
    18256, 
    1, 
    18252, 
    1, 
    18248, 
    1, 
    18245, 
    1, 
    18241, 
    1, 
    18238, 
    1, 
    18234, 
    1, 
    18231, 
    1, 
    18227, 
    1, 
    18223, 
    1, 
    18221, 
    1, 
    18217, 
    1, 
    18213, 
    1, 
    18210, 
    1, 
    18206, 
    1, 
    18203, 
    1, 
    18199, 
    1, 
    18196, 
    1, 
    18192, 
    1, 
    18188, 
    1, 
    18186, 
    1, 
    18182, 
    1, 
    18178, 
    1, 
    18175, 
    1, 
    18171, 
    1, 
    18168, 
    1, 
    18164, 
    1, 
    18161, 
    1, 
    18157, 
    1, 
    18153, 
    1, 
    18151, 
    1, 
    18147, 
    1, 
    18143, 
    1, 
    18140, 
    1, 
    18136, 
    1, 
    18133, 
    1, 
    18129, 
    1, 
    18126, 
    1, 
    18122, 
    1, 
    18118, 
    1, 
    18116, 
    1, 
    18112, 
    1, 
    18108, 
    1, 
    18105, 
    1, 
    18101, 
    1, 
    18098, 
    1, 
    18094, 
    1, 
    18094, 
    1, 
    18092, 
    1, 
    18090, 
    1, 
    18090, 
    1, 
    18088, 
    1, 
    18087, 
    1, 
    18086, 
    1, 
    18084, 
    1, 
    18083, 
    1, 
    18081, 
    1, 
    18081, 
    1, 
    18079, 
    1, 
    18077, 
    1, 
    18077, 
    1, 
    18075, 
    1, 
    18074, 
    1, 
    18073, 
    1, 
    18071, 
    1, 
    18070, 
    1, 
    18068, 
    1, 
    18068, 
    1, 
    18066, 
    1, 
    18064, 
    1, 
    18064, 
    1, 
    18062, 
    1, 
    18061, 
    1, 
    18060, 
    1, 
    18058, 
    1, 
    18057, 
    1, 
    18055, 
    1, 
    18055, 
    1, 
    18053, 
    1, 
    18051, 
    1, 
    18051, 
    1, 
    18049, 
    1, 
    18048, 
    1, 
    18047, 
    1, 
    18045, 
    1, 
    18044, 
    1, 
    18042, 
    1, 
    18042, 
    1, 
    18040, 
    1, 
    18038, 
    1, 
    18038, 
    1, 
    18036, 
    1, 
    18035, 
    1, 
    18034, 
    1, 
    18032, 
    1, 
    18031, 
    1, 
    18029, 
    1, 
    18029, 
    1, 
    18027, 
    1, 
    18025, 
    1, 
    18025, 
    1, 
    18023, 
    1, 
    18022, 
    1, 
    18021, 
    1, 
    18019, 
    1, 
    18018, 
    1, 
    18016, 
    1, 
    18016, 
    1, 
    18014, 
    1, 
    18012, 
    1, 
    18012, 
    1, 
    18010, 
    1, 
    18009, 
    1, 
    18008, 
    1, 
    18006, 
    1, 
    18005, 
    1, 
    18003, 
    1, 
    18003, 
    1, 
    18001, 
    1, 
    17999, 
    1, 
    17999, 
    1, 
    17997, 
    1, 
    17996, 
    1, 
    17995, 
    1, 
    17993, 
    1, 
    17992, 
    1, 
    17990, 
    1, 
    17990, 
    1, 
    17988, 
    1, 
    17986, 
    1, 
    17986, 
    1, 
    17984, 
    1, 
    17983, 
    1, 
    17982, 
    1, 
    17980, 
    1, 
    17979, 
    1, 
    17977, 
    1, 
    17977, 
    1, 
    17975, 
    1, 
    17973, 
    1, 
    17973, 
    1, 
    17971, 
    1, 
    17970, 
    1, 
    17969, 
    1, 
    17967, 
    1, 
    17966, 
    1, 
    17964, 
    1, 
    17964, 
    1, 
    17962, 
    1, 
    17960, 
    1, 
    17960, 
    1, 
    17958, 
    1, 
    17957, 
    1, 
    17956, 
    1, 
    17954, 
    1, 
    17953, 
    1, 
    17951, 
    1, 
    17951, 
    1, 
    17949, 
    1, 
    17947, 
    1, 
    17947, 
    1, 
    17945, 
    1, 
    17944, 
    1, 
    17943, 
    1, 
    17941, 
    1, 
    17940, 
    1, 
    17938, 
    1, 
    17938, 
    1, 
    17936, 
    1, 
    17934, 
    1, 
    17934, 
    1, 
    17932, 
    1, 
    17931, 
    1, 
    17930, 
    1, 
    17928, 
    1, 
    17927, 
    1, 
    17925, 
    1, 
    17925, 
    1, 
    17923, 
    1, 
    17921, 
    1, 
    17921, 
    1, 
    17919, 
    1, 
    17918, 
    1, 
    17917, 
    1, 
    17915, 
    1, 
    17914, 
    1, 
    17912, 
    1, 
    17912, 
    1, 
    17910, 
    1, 
    17908, 
    1, 
    17908, 
    1, 
    17906, 
    1, 
    17905, 
    1, 
    17904, 
    1, 
    17902, 
    1, 
    17901, 
    1, 
    17901, 
    1, 
    17904, 
    1, 
    17907, 
    1, 
    17910, 
    1, 
    17914, 
    1, 
    17917, 
    1, 
    17920, 
    1, 
    17924, 
    1, 
    17927, 
    1, 
    17930, 
    1, 
    17934, 
    1, 
    17937, 
    1, 
    17939, 
    1, 
    17943, 
    1, 
    17946, 
    1, 
    17949, 
    1, 
    17952, 
    1, 
    17956, 
    1, 
    17959, 
    1, 
    17962, 
    1, 
    17966, 
    1, 
    17969, 
    1, 
    17972, 
    1, 
    17975, 
    1, 
    17979, 
    1, 
    17982, 
    1, 
    17985, 
    1, 
    17989, 
    1, 
    17992, 
    1, 
    17995, 
    1, 
    17999, 
    1, 
    18002, 
    1, 
    18005, 
    1, 
    18008, 
    1, 
    18012, 
    1, 
    18015, 
    1, 
    18017, 
    1, 
    18021, 
    1, 
    18024, 
    1, 
    18027, 
    1, 
    18031, 
    1, 
    18034, 
    1, 
    18037, 
    1, 
    18040, 
    1, 
    18044, 
    1, 
    18047, 
    1, 
    18050, 
    1, 
    18054, 
    1, 
    18057, 
    1, 
    18060, 
    1, 
    18064, 
    1, 
    18067, 
    1, 
    18070, 
    1, 
    18073, 
    1, 
    18077, 
    1, 
    18080, 
    1, 
    18083, 
    1, 
    18086, 
    1, 
    18089, 
    1, 
    18092, 
    1, 
    18096, 
    1, 
    18099, 
    1, 
    18102, 
    1, 
    18105, 
    1, 
    18109, 
    1, 
    18112, 
    1, 
    18115, 
    1, 
    18119, 
    1, 
    18122, 
    1, 
    18125, 
    1, 
    18129, 
    1, 
    18132, 
    1, 
    18135, 
    1, 
    18138, 
    1, 
    18140, 
    1, 
    18141, 
    1, 
    18142, 
    1, 
    18144, 
    1, 
    18144, 
    1, 
    18145, 
    1, 
    18147, 
    1, 
    18148, 
    1, 
    18149, 
    1, 
    18150, 
    1, 
    18152, 
    1, 
    18153, 
    1, 
    18153, 
    1, 
    18155, 
    1, 
    18156, 
    1, 
    18157, 
    1, 
    18159, 
    1, 
    18160, 
    1, 
    18161, 
    1, 
    18162, 
    1, 
    18163, 
    1, 
    18164, 
    1, 
    18165, 
    1, 
    18167, 
    1, 
    18168, 
    1, 
    18169, 
    1, 
    18171, 
    1, 
    18172, 
    1, 
    18172, 
    1, 
    18173, 
    1, 
    18175, 
    1, 
    18176, 
    1, 
    18177, 
    1, 
    18179, 
    1, 
    18180, 
    1, 
    18181, 
    1, 
    18182, 
    1, 
    18183, 
    1, 
    18184, 
    1, 
    18185, 
    1, 
    18187, 
    1, 
    18188, 
    1, 
    18189, 
    1, 
    18191, 
    1, 
    18191, 
    1, 
    18192, 
    1, 
    18194, 
    1, 
    18195, 
    1, 
    18196, 
    1, 
    18197, 
    1, 
    18199, 
    1, 
    18200, 
    1, 
    18200, 
    1, 
    18204, 
    1, 
    18208, 
    1, 
    18211, 
    1, 
    18216, 
    1, 
    18220, 
    1, 
    18224, 
    1, 
    18228, 
    1, 
    18232, 
    1, 
    18236, 
    1, 
    18240, 
    1, 
    18245, 
    1, 
    18249, 
    1, 
    18252, 
    1, 
    18257, 
    1, 
    18261, 
    1, 
    18265, 
    1, 
    18269, 
    1, 
    18274, 
    1, 
    18279, 
    1, 
    18283, 
    1, 
    18289, 
    1, 
    18294, 
    1, 
    18298, 
    1, 
    18304, 
    1, 
    18309, 
    1, 
    18313, 
    1, 
    18318, 
    1, 
    18324, 
    1, 
    18328, 
    1, 
    18333, 
    1, 
    18339, 
    1, 
    18343, 
    1, 
    18348, 
    1, 
    18354, 
    1, 
    18358, 
    1, 
    18363, 
    1, 
    18368, 
    1, 
    18372, 
    1, 
    18374, 
    1, 
    18376, 
    1, 
    18380, 
    1, 
    18382, 
    1, 
    18385, 
    1, 
    18388, 
    1, 
    18390, 
    1, 
    18393, 
    1, 
    18395, 
    1, 
    18399, 
    1, 
    18401, 
    1, 
    18403, 
    1, 
    18407, 
    1, 
    18409, 
    1, 
    18412, 
    1, 
    18415, 
    1, 
    18417, 
    1, 
    18420, 
    1, 
    18422, 
    1, 
    18426, 
    1, 
    18430, 
    1, 
    18434, 
    1, 
    18440, 
    1, 
    18445, 
    1, 
    18450, 
    1, 
    18455, 
    1, 
    18459, 
    1, 
    18465, 
    1, 
    18469, 
    1, 
    18474, 
    1, 
    18479, 
    1, 
    18484, 
    1, 
    18490, 
    1, 
    18496, 
    1, 
    18503, 
    1, 
    18509, 
    1, 
    18516, 
    1, 
    18521, 
    1, 
    18528, 
    1, 
    18534, 
    1, 
    18541, 
    1, 
    18547, 
    1, 
    18553, 
    1, 
    18560, 
    1, 
    18566, 
    1, 
    18573, 
    1, 
    18578, 
    1, 
    18585, 
    1, 
    18591, 
    1, 
    18598, 
    1, 
    18604, 
    1, 
    18610, 
    1, 
    18617, 
    1, 
    18623, 
    1, 
    18630, 
    1, 
    18635, 
    1, 
    18642, 
    1, 
    18648, 
    1, 
    18655, 
    1, 
    18661, 
    1, 
    18667, 
    1, 
    18674, 
    1, 
    18681, 
    1, 
    18689, 
    1, 
    18697, 
    1, 
    18705, 
    1, 
    18712, 
    1, 
    18721, 
    1, 
    18729, 
    1, 
    18737, 
    1, 
    18745, 
    1, 
    18753, 
    1, 
    18761, 
    1, 
    18768, 
    1, 
    18777, 
    1, 
    18784, 
    1, 
    18793, 
    1, 
    18800, 
    1, 
    18808, 
    1, 
    18817, 
    1, 
    18824, 
    1, 
    18833, 
    1, 
    18840, 
    1, 
    18849, 
    1, 
    18856, 
    1, 
    18864, 
    1, 
    18872, 
    1, 
    18880, 
    1, 
    18889, 
    1, 
    18896, 
    1, 
    18905, 
    1, 
    18912, 
    1, 
    18920, 
    1, 
    18928, 
    1, 
    18936, 
    1, 
    18944, 
    1, 
    18952, 
    1, 
    18960, 
    1, 
    18968, 
    1, 
    18976, 
    1, 
    18984, 
    1, 
    18992, 
    1, 
    19000, 
    1, 
    19008, 
    1, 
    19016, 
    1, 
    19024, 
    1, 
    19032, 
    1, 
    19040, 
    1, 
    19048, 
    1, 
    19056, 
    1, 
    19064, 
    1, 
    19071, 
    1, 
    19080, 
    1, 
    19087, 
    1, 
    19096, 
    1, 
    19104, 
    1, 
    19112, 
    1, 
    19120, 
    1, 
    19127, 
    1, 
    19136, 
    1, 
    19143, 
    1, 
    19152, 
    1, 
    19159, 
    1, 
    19168, 
    1, 
    19176, 
    1, 
    19183, 
    1, 
    19192, 
    1, 
    19199, 
    1, 
    19208, 
    1, 
    19215, 
    1, 
    19224, 
    1, 
    19231, 
    1, 
    19239, 
    1, 
    19248, 
    1, 
    19255, 
    1, 
    19264, 
    1, 
    19271, 
    1, 
    19279, 
    1, 
    19287, 
    1, 
    19295, 
    1, 
    19303, 
    1, 
    19311, 
    1, 
    19320, 
    1, 
    19327, 
    1, 
    19336, 
    1, 
    19343, 
    1, 
    19351, 
    1, 
    19359, 
    1, 
    19367, 
    1, 
    19375, 
    1, 
    19383, 
    1, 
    19391, 
    1, 
    19399, 
    1, 
    19407, 
    1, 
    19415, 
    1, 
    19423, 
    1, 
    19431, 
    1, 
    19439, 
    1, 
    19446, 
    1, 
    19455, 
    1, 
    19463, 
    1, 
    19471, 
    1, 
    19479, 
    1, 
    19487, 
    1, 
    19495, 
    1, 
    19502, 
    1, 
    19511, 
    1, 
    19518, 
    1, 
    19527, 
    1, 
    19534, 
    1, 
    19543, 
    1, 
    19551, 
    1, 
    19558, 
    1, 
    19567, 
    1, 
    19574, 
    1, 
    19583, 
    1, 
    19590, 
    1, 
    19598, 
    1, 
    19606, 
    1, 
    19614, 
    1, 
    19623, 
    1, 
    19630, 
    1, 
    19639, 
    1, 
    19646, 
    1, 
    19654, 
    1, 
    19662, 
    1, 
    19670, 
    1, 
    19678, 
    1, 
    19686, 
    1, 
    19695, 
    1, 
    19702, 
    1, 
    19710, 
    1, 
    19718, 
    1, 
    19726, 
    1, 
    19734, 
    1, 
    19742, 
    1, 
    19750, 
    1, 
    19758, 
    1, 
    19766, 
    1, 
    19774, 
    1, 
    19782, 
    1, 
    19790, 
    1, 
    19798, 
    1, 
    19806, 
    1, 
    19814, 
    1, 
    19821, 
    1, 
    19830, 
    1, 
    19838, 
    1, 
    19846, 
    1, 
    19854, 
    1, 
    19862, 
    1, 
    19870, 
    1, 
    19877, 
    1, 
    19886, 
    1, 
    19893, 
    1, 
    19902, 
    1, 
    19910, 
    1, 
    19917, 
    1, 
    19926, 
    1, 
    19933, 
    1, 
    19942, 
    1, 
    19949, 
    1, 
    19958, 
    1, 
    19965, 
    1, 
    19973, 
    1, 
    19982, 
    1, 
    19989, 
    1, 
    19998, 
    1, 
    20005, 
    1, 
    20014, 
    1, 
    20021, 
    1, 
    20029, 
    1, 
    20037, 
    1, 
    20045, 
    1, 
    20054, 
    1, 
    20061, 
    1, 
    20070, 
    1, 
    20077, 
    1, 
    20085, 
    1, 
    20093, 
    1, 
    20101, 
    1, 
    20109, 
    1, 
    20117, 
    1, 
    20126, 
    1, 
    20133, 
    1, 
    20141, 
    1, 
    20149, 
    1, 
    20157, 
    1, 
    20165, 
    1, 
    20173, 
    1, 
    20181, 
    1, 
    20189, 
    1, 
    20197, 
    1, 
    20205, 
    1, 
    20213, 
    1, 
    20221, 
    1, 
    20229, 
    1, 
    20236, 
    1, 
    20245, 
    1, 
    20252, 
    1, 
    20261, 
    1, 
    20268, 
    1, 
    20277, 
    1, 
    20285, 
    1, 
    20292, 
    1, 
    20301, 
    1, 
    20308, 
    1, 
    20317, 
    1, 
    20324, 
    1, 
    20333, 
    1, 
    20340, 
    1, 
    20348, 
    1, 
    20357, 
    1, 
    20364, 
    1, 
    20373, 
    1, 
    20380, 
    1, 
    20389, 
    1, 
    20396, 
    1, 
    20404, 
    1, 
    20412, 
    1, 
    20420, 
    1, 
    20429, 
    1, 
    20436, 
    1, 
    20445, 
    1, 
    20452, 
    1, 
    20460, 
    1, 
    20468, 
    1, 
    20476, 
    1, 
    20484, 
    1, 
    20492, 
    1, 
    20501, 
    1, 
    20508, 
    1, 
    20516, 
    1, 
    20524, 
    1, 
    20532, 
    1, 
    20540, 
    1, 
    20548, 
    1, 
    20555, 
    1, 
    20564, 
    1, 
    20572, 
    1, 
    20580, 
    1, 
    20588, 
    1, 
    20596, 
    1, 
    20604, 
    1, 
    20611, 
    1, 
    20627, 
    1, 
    20676, 
    1, 
    20726, 
    1, 
    20774, 
    1, 
    20823, 
    1, 
    20872, 
    1, 
    20922, 
    1, 
    20970, 
    1, 
    21019, 
    1, 
    21069, 
    1, 
    21118, 
    1, 
    21166, 
    1, 
    21216, 
    1, 
    21265, 
    1, 
    21314, 
    1, 
    21362, 
    1, 
    21412, 
    1, 
    21461, 
    1, 
    21510, 
    1, 
    21558, 1 ;
}
